library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

--library UNISIM;
--use UNISIM.VComponents.all;

entity OUTPUT_LAYER is
Generic (WIDTH : positive := 32);
Port (
     CLK     :  in std_logic;
     RESET   :  in std_logic;
     SET_CNT :  in std_logic;
     DIN0    :  in std_logic_vector(WIDTH-1 downto 0);
     DIN1    :  in std_logic_vector(WIDTH-1 downto 0);
     DIN2    :  in std_logic_vector(WIDTH-1 downto 0);
     DIN3    :  in std_logic_vector(WIDTH-1 downto 0);
     DIN4    :  in std_logic_vector(WIDTH-1 downto 0);
     DIN5    :  in std_logic_vector(WIDTH-1 downto 0);
     DIN6    :  in std_logic_vector(WIDTH-1 downto 0);
     DIN7    :  in std_logic_vector(WIDTH-1 downto 0);
     DIN8    :  in std_logic_vector(WIDTH-1 downto 0);
     DIN9    :  in std_logic_vector(WIDTH-1 downto 0);
     DIN10   :  in std_logic_vector(WIDTH-1 downto 0);
     DIN11   :  in std_logic_vector(WIDTH-1 downto 0);
     DIN12   :  in std_logic_vector(WIDTH-1 downto 0);
     DIN13   :  in std_logic_vector(WIDTH-1 downto 0);
     DIN14   :  in std_logic_vector(WIDTH-1 downto 0);
     DIN15   :  in std_logic_vector(WIDTH-1 downto 0);
     DIN16   :  in std_logic_vector(WIDTH-1 downto 0);
     DIN17   :  in std_logic_vector(WIDTH-1 downto 0);
     DIN18   :  in std_logic_vector(WIDTH-1 downto 0);
     DIN19   :  in std_logic_vector(WIDTH-1 downto 0);
     DIN20   :  in std_logic_vector(WIDTH-1 downto 0);
     DIN21   :  in std_logic_vector(WIDTH-1 downto 0);
     DIN22   :  in std_logic_vector(WIDTH-1 downto 0);
     DIN23   :  in std_logic_vector(WIDTH-1 downto 0);
     DIN24   :  in std_logic_vector(WIDTH-1 downto 0);
     DIN25   :  in std_logic_vector(WIDTH-1 downto 0);
     DIN26   :  in std_logic_vector(WIDTH-1 downto 0);
     DIN27   :  in std_logic_vector(WIDTH-1 downto 0);
     DIN28   :  in std_logic_vector(WIDTH-1 downto 0);
     DIN29   :  in std_logic_vector(WIDTH-1 downto 0);
     DOUT0   :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
     DOUT1   :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
     DOUT2   :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
     DOUT3   :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
     DOUT4   :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
     DOUT5   :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
     DOUT6   :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
     DOUT7   :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
     DOUT8   :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
     DOUT9   :  out std_logic_vector(WIDTH+WIDTH-1 downto 0)
);
end OUTPUT_LAYER;

architecture Structural of OUTPUT_LAYER is

component OUTPUT_VECTOR_MULTIPLIER
Generic(WIDTH : positive := 32;
        POWER : positive := 5);
Port (
    CLK         :  in  std_logic;
    RESET       :  in  std_logic;
    SET         :  in  std_logic;
    DIN0        :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN1        :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN2        :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN3        :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN4        :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN5        :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN6        :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN7        :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN8        :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN9        :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN10       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN11       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN12       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN13       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN14       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN15       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN16       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN17       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN18       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN19       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN20       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN21       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN22       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN23       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN24       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN25       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN26       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN27       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN28       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN29       :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM0_DATA   :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM1_DATA   :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM2_DATA   :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM3_DATA   :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM4_DATA   :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM5_DATA   :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM6_DATA   :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM7_DATA   :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM8_DATA   :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM9_DATA   :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM10_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM11_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM12_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM13_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM14_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM15_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM16_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM17_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM18_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM19_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM20_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM21_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM22_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM23_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM24_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM25_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM26_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM27_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM28_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM29_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ADDR0       :  out std_logic_vector(POWER-1 downto 0);
    ADDR1       :  out std_logic_vector(POWER-1 downto 0);
    ADDR2       :  out std_logic_vector(POWER-1 downto 0);
    ADDR3       :  out std_logic_vector(POWER-1 downto 0);
    ADDR4       :  out std_logic_vector(POWER-1 downto 0);
    ADDR5       :  out std_logic_vector(POWER-1 downto 0);
    ADDR6       :  out std_logic_vector(POWER-1 downto 0);
    ADDR7       :  out std_logic_vector(POWER-1 downto 0);
    ADDR8       :  out std_logic_vector(POWER-1 downto 0);
    ADDR9       :  out std_logic_vector(POWER-1 downto 0);
    ADDR10      :  out std_logic_vector(POWER-1 downto 0);
    ADDR11      :  out std_logic_vector(POWER-1 downto 0);
    ADDR12      :  out std_logic_vector(POWER-1 downto 0);
    ADDR13      :  out std_logic_vector(POWER-1 downto 0);
    ADDR14      :  out std_logic_vector(POWER-1 downto 0);
    ADDR15      :  out std_logic_vector(POWER-1 downto 0);
    ADDR16      :  out std_logic_vector(POWER-1 downto 0);
    ADDR17      :  out std_logic_vector(POWER-1 downto 0);
    ADDR18      :  out std_logic_vector(POWER-1 downto 0);
    ADDR19      :  out std_logic_vector(POWER-1 downto 0);
    ADDR20      :  out std_logic_vector(POWER-1 downto 0);
    ADDR21      :  out std_logic_vector(POWER-1 downto 0);
    ADDR22      :  out std_logic_vector(POWER-1 downto 0);
    ADDR23      :  out std_logic_vector(POWER-1 downto 0);
    ADDR24      :  out std_logic_vector(POWER-1 downto 0);
    ADDR25      :  out std_logic_vector(POWER-1 downto 0);
    ADDR26      :  out std_logic_vector(POWER-1 downto 0);
    ADDR27      :  out std_logic_vector(POWER-1 downto 0);
    ADDR28      :  out std_logic_vector(POWER-1 downto 0);
    ADDR29      :  out std_logic_vector(POWER-1 downto 0);
    DOUT        :  out std_logic_vector(WIDTH+WIDTH-1 downto 0)
);
end component;

component OUTPUT_WEIGHT_ROM
Generic ( WIDTH : positive := 32;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR26 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR27 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR28 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR29 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0);
    DATA26 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA27 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA28 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA29 :    out std_logic_vector(WIDTH-1 downto 0)
);
end component;

component OUTPUT_BIAS_ROM 
Generic ( WIDTH : positive := 64;
          POWER : positive := 4); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0)
);
end component;

component ADDER
Generic ( WIDTH : positive := 32);
Port (
    A    :  in  std_logic_vector(WIDTH-1 downto 0);
    B    :  in  std_logic_vector(WIDTH-1 downto 0);
    S    :  out std_logic_vector(WIDTH-1 downto 0);
    COUT :  out std_logic;
    OV   :  out std_logic
);
end component;

component RELU_MUX
Generic( WIDTH : positive := 32);
Port (
    DIN  :  in  std_logic_vector(WIDTH-1 downto 0);
    DOUT :  out std_logic_vector(WIDTH-1 downto 0)
);
end component;

signal DIN0_SIG, DIN1_SIG, DIN2_SIG, DIN3_SIG, DIN4_SIG, DIN5_SIG, DIN6_SIG, DIN7_SIG, DIN8_SIG,
       DIN9_SIG, DIN10_SIG, DIN11_SIG, DIN12_SIG, DIN13_SIG, DIN14_SIG, DIN15_SIG, DIN16_SIG, DIN17_SIG,
       DIN18_SIG, DIN19_SIG, DIN20_SIG, DIN21_SIG, DIN22_SIG, DIN23_SIG, DIN24_SIG, DIN25_SIG, DIN26_SIG,
       DIN27_SIG, DIN28_SIG, DIN29_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM0_DATA0_SIG,  ROM0_DATA1_SIG,  ROM0_DATA2_SIG,  ROM0_DATA3_SIG,  ROM0_DATA4_SIG,
       ROM0_DATA5_SIG,  ROM0_DATA6_SIG,  ROM0_DATA7_SIG,  ROM0_DATA8_SIG,  ROM0_DATA9_SIG,
       ROM0_DATA10_SIG, ROM0_DATA11_SIG, ROM0_DATA12_SIG, ROM0_DATA13_SIG, ROM0_DATA14_SIG,
       ROM0_DATA15_SIG, ROM0_DATA16_SIG, ROM0_DATA17_SIG, ROM0_DATA18_SIG, ROM0_DATA19_SIG,
       ROM0_DATA20_SIG, ROM0_DATA21_SIG, ROM0_DATA22_SIG, ROM0_DATA23_SIG, ROM0_DATA24_SIG,
       ROM0_DATA25_SIG, ROM0_DATA26_SIG, ROM0_DATA27_SIG, ROM0_DATA28_SIG,  ROM0_DATA29_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM1_DATA0_SIG,  ROM1_DATA1_SIG,  ROM1_DATA2_SIG,  ROM1_DATA3_SIG,  ROM1_DATA4_SIG,
       ROM1_DATA5_SIG,  ROM1_DATA6_SIG,  ROM1_DATA7_SIG,  ROM1_DATA8_SIG,  ROM1_DATA9_SIG,
       ROM1_DATA10_SIG, ROM1_DATA11_SIG, ROM1_DATA12_SIG, ROM1_DATA13_SIG, ROM1_DATA14_SIG,
       ROM1_DATA15_SIG, ROM1_DATA16_SIG, ROM1_DATA17_SIG, ROM1_DATA18_SIG, ROM1_DATA19_SIG,
       ROM1_DATA20_SIG, ROM1_DATA21_SIG, ROM1_DATA22_SIG, ROM1_DATA23_SIG, ROM1_DATA24_SIG,
       ROM1_DATA25_SIG, ROM1_DATA26_SIG, ROM1_DATA27_SIG, ROM1_DATA28_SIG,  ROM1_DATA29_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM2_DATA0_SIG,  ROM2_DATA1_SIG,  ROM2_DATA2_SIG,  ROM2_DATA3_SIG,  ROM2_DATA4_SIG,
       ROM2_DATA5_SIG,  ROM2_DATA6_SIG,  ROM2_DATA7_SIG,  ROM2_DATA8_SIG,  ROM2_DATA9_SIG,
       ROM2_DATA10_SIG, ROM2_DATA11_SIG, ROM2_DATA12_SIG, ROM2_DATA13_SIG, ROM2_DATA14_SIG,
       ROM2_DATA15_SIG, ROM2_DATA16_SIG, ROM2_DATA17_SIG, ROM2_DATA18_SIG, ROM2_DATA19_SIG,
       ROM2_DATA20_SIG, ROM2_DATA21_SIG, ROM2_DATA22_SIG, ROM2_DATA23_SIG, ROM2_DATA24_SIG,
       ROM2_DATA25_SIG, ROM2_DATA26_SIG, ROM2_DATA27_SIG, ROM2_DATA28_SIG,  ROM2_DATA29_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM3_DATA0_SIG,  ROM3_DATA1_SIG,  ROM3_DATA2_SIG,  ROM3_DATA3_SIG,  ROM3_DATA4_SIG,
       ROM3_DATA5_SIG,  ROM3_DATA6_SIG,  ROM3_DATA7_SIG,  ROM3_DATA8_SIG,  ROM3_DATA9_SIG,
       ROM3_DATA10_SIG, ROM3_DATA11_SIG, ROM3_DATA12_SIG, ROM3_DATA13_SIG, ROM3_DATA14_SIG,
       ROM3_DATA15_SIG, ROM3_DATA16_SIG, ROM3_DATA17_SIG, ROM3_DATA18_SIG, ROM3_DATA19_SIG,
       ROM3_DATA20_SIG, ROM3_DATA21_SIG, ROM3_DATA22_SIG, ROM3_DATA23_SIG, ROM3_DATA24_SIG,
       ROM3_DATA25_SIG, ROM3_DATA26_SIG, ROM3_DATA27_SIG, ROM3_DATA28_SIG,  ROM3_DATA29_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM4_DATA0_SIG,  ROM4_DATA1_SIG,  ROM4_DATA2_SIG,  ROM4_DATA3_SIG,  ROM4_DATA4_SIG,
       ROM4_DATA5_SIG,  ROM4_DATA6_SIG,  ROM4_DATA7_SIG,  ROM4_DATA8_SIG,  ROM4_DATA9_SIG,
       ROM4_DATA10_SIG, ROM4_DATA11_SIG, ROM4_DATA12_SIG, ROM4_DATA13_SIG, ROM4_DATA14_SIG,
       ROM4_DATA15_SIG, ROM4_DATA16_SIG, ROM4_DATA17_SIG, ROM4_DATA18_SIG, ROM4_DATA19_SIG,
       ROM4_DATA20_SIG, ROM4_DATA21_SIG, ROM4_DATA22_SIG, ROM4_DATA23_SIG, ROM4_DATA24_SIG,
       ROM4_DATA25_SIG, ROM4_DATA26_SIG, ROM4_DATA27_SIG, ROM4_DATA28_SIG,  ROM4_DATA29_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM5_DATA0_SIG,  ROM5_DATA1_SIG,  ROM5_DATA2_SIG,  ROM5_DATA3_SIG,  ROM5_DATA4_SIG,
       ROM5_DATA5_SIG,  ROM5_DATA6_SIG,  ROM5_DATA7_SIG,  ROM5_DATA8_SIG,  ROM5_DATA9_SIG,
       ROM5_DATA10_SIG, ROM5_DATA11_SIG, ROM5_DATA12_SIG, ROM5_DATA13_SIG, ROM5_DATA14_SIG,
       ROM5_DATA15_SIG, ROM5_DATA16_SIG, ROM5_DATA17_SIG, ROM5_DATA18_SIG, ROM5_DATA19_SIG,
       ROM5_DATA20_SIG, ROM5_DATA21_SIG, ROM5_DATA22_SIG, ROM5_DATA23_SIG, ROM5_DATA24_SIG,
       ROM5_DATA25_SIG, ROM5_DATA26_SIG, ROM5_DATA27_SIG, ROM5_DATA28_SIG,  ROM5_DATA29_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM6_DATA0_SIG,  ROM6_DATA1_SIG,  ROM6_DATA2_SIG,  ROM6_DATA3_SIG,  ROM6_DATA4_SIG,
       ROM6_DATA5_SIG,  ROM6_DATA6_SIG,  ROM6_DATA7_SIG,  ROM6_DATA8_SIG,  ROM6_DATA9_SIG,
       ROM6_DATA10_SIG, ROM6_DATA11_SIG, ROM6_DATA12_SIG, ROM6_DATA13_SIG, ROM6_DATA14_SIG,
       ROM6_DATA15_SIG, ROM6_DATA16_SIG, ROM6_DATA17_SIG, ROM6_DATA18_SIG, ROM6_DATA19_SIG,
       ROM6_DATA20_SIG, ROM6_DATA21_SIG, ROM6_DATA22_SIG, ROM6_DATA23_SIG, ROM6_DATA24_SIG,
       ROM6_DATA25_SIG, ROM6_DATA26_SIG, ROM6_DATA27_SIG, ROM6_DATA28_SIG,  ROM6_DATA29_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM7_DATA0_SIG,  ROM7_DATA1_SIG,  ROM7_DATA2_SIG,  ROM7_DATA3_SIG,  ROM7_DATA4_SIG,
       ROM7_DATA5_SIG,  ROM7_DATA6_SIG,  ROM7_DATA7_SIG,  ROM7_DATA8_SIG,  ROM7_DATA9_SIG,
       ROM7_DATA10_SIG, ROM7_DATA11_SIG, ROM7_DATA12_SIG, ROM7_DATA13_SIG, ROM7_DATA14_SIG,
       ROM7_DATA15_SIG, ROM7_DATA16_SIG, ROM7_DATA17_SIG, ROM7_DATA18_SIG, ROM7_DATA19_SIG,
       ROM7_DATA20_SIG, ROM7_DATA21_SIG, ROM7_DATA22_SIG, ROM7_DATA23_SIG, ROM7_DATA24_SIG,
       ROM7_DATA25_SIG, ROM7_DATA26_SIG, ROM7_DATA27_SIG, ROM7_DATA28_SIG,  ROM7_DATA29_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM8_DATA0_SIG,  ROM8_DATA1_SIG,  ROM8_DATA2_SIG,  ROM8_DATA3_SIG,  ROM8_DATA4_SIG,
       ROM8_DATA5_SIG,  ROM8_DATA6_SIG,  ROM8_DATA7_SIG,  ROM8_DATA8_SIG,  ROM8_DATA9_SIG,
       ROM8_DATA10_SIG, ROM8_DATA11_SIG, ROM8_DATA12_SIG, ROM8_DATA13_SIG, ROM8_DATA14_SIG,
       ROM8_DATA15_SIG, ROM8_DATA16_SIG, ROM8_DATA17_SIG, ROM8_DATA18_SIG, ROM8_DATA19_SIG,
       ROM8_DATA20_SIG, ROM8_DATA21_SIG, ROM8_DATA22_SIG, ROM8_DATA23_SIG, ROM8_DATA24_SIG,
       ROM8_DATA25_SIG, ROM8_DATA26_SIG, ROM8_DATA27_SIG, ROM8_DATA28_SIG,  ROM8_DATA29_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM9_DATA0_SIG,  ROM9_DATA1_SIG,  ROM9_DATA2_SIG,  ROM9_DATA3_SIG,  ROM9_DATA4_SIG,
       ROM9_DATA5_SIG,  ROM9_DATA6_SIG,  ROM9_DATA7_SIG,  ROM9_DATA8_SIG,  ROM9_DATA9_SIG,
       ROM9_DATA10_SIG, ROM9_DATA11_SIG, ROM9_DATA12_SIG, ROM9_DATA13_SIG, ROM9_DATA14_SIG,
       ROM9_DATA15_SIG, ROM9_DATA16_SIG, ROM9_DATA17_SIG, ROM9_DATA18_SIG, ROM9_DATA19_SIG,
       ROM9_DATA20_SIG, ROM9_DATA21_SIG, ROM9_DATA22_SIG, ROM9_DATA23_SIG, ROM9_DATA24_SIG,
       ROM9_DATA25_SIG, ROM9_DATA26_SIG, ROM9_DATA27_SIG, ROM9_DATA28_SIG,  ROM9_DATA29_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ADDR0_0_SIG,  ADDR0_1_SIG,  ADDR0_2_SIG,  ADDR0_3_SIG,  ADDR0_4_SIG,  ADDR0_5_SIG,
       ADDR0_6_SIG,  ADDR0_7_SIG,  ADDR0_8_SIG,  ADDR0_9_SIG,  ADDR0_10_SIG, ADDR0_11_SIG,
       ADDR0_12_SIG, ADDR0_13_SIG, ADDR0_14_SIG, ADDR0_15_SIG, ADDR0_16_SIG, ADDR0_17_SIG,
       ADDR0_18_SIG, ADDR0_19_SIG, ADDR0_20_SIG, ADDR0_21_SIG, ADDR0_22_SIG, ADDR0_23_SIG,
       ADDR0_24_SIG, ADDR0_25_SIG, ADDR0_26_SIG, ADDR0_27_SIG, ADDR0_28_SIG, ADDR0_29_SIG : std_logic_vector(4 downto 0) := (others => '0');
signal ADDR1_0_SIG,  ADDR1_1_SIG,  ADDR1_2_SIG,  ADDR1_3_SIG,  ADDR1_4_SIG,  ADDR1_5_SIG,
       ADDR1_6_SIG,  ADDR1_7_SIG,  ADDR1_8_SIG,  ADDR1_9_SIG,  ADDR1_10_SIG, ADDR1_11_SIG,
       ADDR1_12_SIG, ADDR1_13_SIG, ADDR1_14_SIG, ADDR1_15_SIG, ADDR1_16_SIG, ADDR1_17_SIG,
       ADDR1_18_SIG, ADDR1_19_SIG, ADDR1_20_SIG, ADDR1_21_SIG, ADDR1_22_SIG, ADDR1_23_SIG,
       ADDR1_24_SIG, ADDR1_25_SIG, ADDR1_26_SIG, ADDR1_27_SIG, ADDR1_28_SIG, ADDR1_29_SIG : std_logic_vector(4 downto 0) := (others => '0');
signal ADDR2_0_SIG,  ADDR2_1_SIG,  ADDR2_2_SIG,  ADDR2_3_SIG,  ADDR2_4_SIG,  ADDR2_5_SIG,
       ADDR2_6_SIG,  ADDR2_7_SIG,  ADDR2_8_SIG,  ADDR2_9_SIG,  ADDR2_10_SIG, ADDR2_11_SIG,
       ADDR2_12_SIG, ADDR2_13_SIG, ADDR2_14_SIG, ADDR2_15_SIG, ADDR2_16_SIG, ADDR2_17_SIG,
       ADDR2_18_SIG, ADDR2_19_SIG, ADDR2_20_SIG, ADDR2_21_SIG, ADDR2_22_SIG, ADDR2_23_SIG,
       ADDR2_24_SIG, ADDR2_25_SIG, ADDR2_26_SIG, ADDR2_27_SIG, ADDR2_28_SIG, ADDR2_29_SIG : std_logic_vector(4 downto 0) := (others => '0');
signal ADDR3_0_SIG,  ADDR3_1_SIG,  ADDR3_2_SIG,  ADDR3_3_SIG,  ADDR3_4_SIG,  ADDR3_5_SIG,
       ADDR3_6_SIG,  ADDR3_7_SIG,  ADDR3_8_SIG,  ADDR3_9_SIG,  ADDR3_10_SIG, ADDR3_11_SIG,
       ADDR3_12_SIG, ADDR3_13_SIG, ADDR3_14_SIG, ADDR3_15_SIG, ADDR3_16_SIG, ADDR3_17_SIG,
       ADDR3_18_SIG, ADDR3_19_SIG, ADDR3_20_SIG, ADDR3_21_SIG, ADDR3_22_SIG, ADDR3_23_SIG,
       ADDR3_24_SIG, ADDR3_25_SIG, ADDR3_26_SIG, ADDR3_27_SIG, ADDR3_28_SIG, ADDR3_29_SIG : std_logic_vector(4 downto 0) := (others => '0');
signal ADDR4_0_SIG,  ADDR4_1_SIG,  ADDR4_2_SIG,  ADDR4_3_SIG,  ADDR4_4_SIG,  ADDR4_5_SIG,
       ADDR4_6_SIG,  ADDR4_7_SIG,  ADDR4_8_SIG,  ADDR4_9_SIG,  ADDR4_10_SIG, ADDR4_11_SIG,
       ADDR4_12_SIG, ADDR4_13_SIG, ADDR4_14_SIG, ADDR4_15_SIG, ADDR4_16_SIG, ADDR4_17_SIG,
       ADDR4_18_SIG, ADDR4_19_SIG, ADDR4_20_SIG, ADDR4_21_SIG, ADDR4_22_SIG, ADDR4_23_SIG,
       ADDR4_24_SIG, ADDR4_25_SIG, ADDR4_26_SIG, ADDR4_27_SIG, ADDR4_28_SIG, ADDR4_29_SIG : std_logic_vector(4 downto 0) := (others => '0');
signal ADDR5_0_SIG,  ADDR5_1_SIG,  ADDR5_2_SIG,  ADDR5_3_SIG,  ADDR5_4_SIG,  ADDR5_5_SIG,
       ADDR5_6_SIG,  ADDR5_7_SIG,  ADDR5_8_SIG,  ADDR5_9_SIG,  ADDR5_10_SIG, ADDR5_11_SIG,
       ADDR5_12_SIG, ADDR5_13_SIG, ADDR5_14_SIG, ADDR5_15_SIG, ADDR5_16_SIG, ADDR5_17_SIG,
       ADDR5_18_SIG, ADDR5_19_SIG, ADDR5_20_SIG, ADDR5_21_SIG, ADDR5_22_SIG, ADDR5_23_SIG,
       ADDR5_24_SIG, ADDR5_25_SIG, ADDR5_26_SIG, ADDR5_27_SIG, ADDR5_28_SIG, ADDR5_29_SIG : std_logic_vector(4 downto 0) := (others => '0');
signal ADDR6_0_SIG,  ADDR6_1_SIG,  ADDR6_2_SIG,  ADDR6_3_SIG,  ADDR6_4_SIG,  ADDR6_5_SIG,
       ADDR6_6_SIG,  ADDR6_7_SIG,  ADDR6_8_SIG,  ADDR6_9_SIG,  ADDR6_10_SIG, ADDR6_11_SIG,
       ADDR6_12_SIG, ADDR6_13_SIG, ADDR6_14_SIG, ADDR6_15_SIG, ADDR6_16_SIG, ADDR6_17_SIG,
       ADDR6_18_SIG, ADDR6_19_SIG, ADDR6_20_SIG, ADDR6_21_SIG, ADDR6_22_SIG, ADDR6_23_SIG,
       ADDR6_24_SIG, ADDR6_25_SIG, ADDR6_26_SIG, ADDR6_27_SIG, ADDR6_28_SIG, ADDR6_29_SIG : std_logic_vector(4 downto 0) := (others => '0');
signal ADDR7_0_SIG,  ADDR7_1_SIG,  ADDR7_2_SIG,  ADDR7_3_SIG,  ADDR7_4_SIG,  ADDR7_5_SIG,
       ADDR7_6_SIG,  ADDR7_7_SIG,  ADDR7_8_SIG,  ADDR7_9_SIG,  ADDR7_10_SIG, ADDR7_11_SIG,
       ADDR7_12_SIG, ADDR7_13_SIG, ADDR7_14_SIG, ADDR7_15_SIG, ADDR7_16_SIG, ADDR7_17_SIG,
       ADDR7_18_SIG, ADDR7_19_SIG, ADDR7_20_SIG, ADDR7_21_SIG, ADDR7_22_SIG, ADDR7_23_SIG,
       ADDR7_24_SIG, ADDR7_25_SIG, ADDR7_26_SIG, ADDR7_27_SIG, ADDR7_28_SIG, ADDR7_29_SIG : std_logic_vector(4 downto 0) := (others => '0');
signal ADDR8_0_SIG,  ADDR8_1_SIG,  ADDR8_2_SIG,  ADDR8_3_SIG,  ADDR8_4_SIG,  ADDR8_5_SIG,
       ADDR8_6_SIG,  ADDR8_7_SIG,  ADDR8_8_SIG,  ADDR8_9_SIG,  ADDR8_10_SIG, ADDR8_11_SIG,
       ADDR8_12_SIG, ADDR8_13_SIG, ADDR8_14_SIG, ADDR8_15_SIG, ADDR8_16_SIG, ADDR8_17_SIG,
       ADDR8_18_SIG, ADDR8_19_SIG, ADDR8_20_SIG, ADDR8_21_SIG, ADDR8_22_SIG, ADDR8_23_SIG,
       ADDR8_24_SIG, ADDR8_25_SIG, ADDR8_26_SIG, ADDR8_27_SIG, ADDR8_28_SIG, ADDR8_29_SIG : std_logic_vector(4 downto 0) := (others => '0');
signal ADDR9_0_SIG,  ADDR9_1_SIG,  ADDR9_2_SIG,  ADDR9_3_SIG,  ADDR9_4_SIG,  ADDR9_5_SIG,
       ADDR9_6_SIG,  ADDR9_7_SIG,  ADDR9_8_SIG,  ADDR9_9_SIG,  ADDR9_10_SIG, ADDR9_11_SIG,
       ADDR9_12_SIG, ADDR9_13_SIG, ADDR9_14_SIG, ADDR9_15_SIG, ADDR9_16_SIG, ADDR9_17_SIG,
       ADDR9_18_SIG, ADDR9_19_SIG, ADDR9_20_SIG, ADDR9_21_SIG, ADDR9_22_SIG, ADDR9_23_SIG,
       ADDR9_24_SIG, ADDR9_25_SIG, ADDR9_26_SIG, ADDR9_27_SIG, ADDR9_28_SIG, ADDR9_29_SIG : std_logic_vector(4 downto 0) := (others => '0');
signal O_VM0_OUT_SIG, O_VM1_OUT_SIG, O_VM2_OUT_SIG, O_VM3_OUT_SIG, O_VM4_OUT_SIG,
       O_VM5_OUT_SIG, O_VM6_OUT_SIG, O_VM7_OUT_SIG, O_VM8_OUT_SIG, O_VM9_OUT_SIG : std_logic_vector(WIDTH+WIDTH-1 downto 0) := (others => '0');
signal ADDER0_OUT_SIG, ADDER1_OUT_SIG, ADDER2_OUT_SIG, ADDER3_OUT_SIG, ADDER4_OUT_SIG,
       ADDER5_OUT_SIG, ADDER6_OUT_SIG, ADDER7_OUT_SIG, ADDER8_OUT_SIG, ADDER9_OUT_SIG : std_logic_vector(WIDTH+WIDTH-1 downto 0) := (others => '0');
signal SET_O_VM : std_logic := '0';
signal BIAS_ADDR0_SIG : std_logic_vector(3 downto 0) := "0000";
signal BIAS_ADDR1_SIG : std_logic_vector(3 downto 0) := "0001";
signal BIAS_ADDR2_SIG : std_logic_vector(3 downto 0) := "0010";
signal BIAS_ADDR3_SIG : std_logic_vector(3 downto 0) := "0011";
signal BIAS_ADDR4_SIG : std_logic_vector(3 downto 0) := "0100";
signal BIAS_ADDR5_SIG : std_logic_vector(3 downto 0) := "0101";
signal BIAS_ADDR6_SIG : std_logic_vector(3 downto 0) := "0110";
signal BIAS_ADDR7_SIG : std_logic_vector(3 downto 0) := "0111";
signal BIAS_ADDR8_SIG : std_logic_vector(3 downto 0) := "1000";
signal BIAS_ADDR9_SIG : std_logic_vector(3 downto 0) := "1001";
signal BIAS0_SIG, BIAS1_SIG, BIAS2_SIG, BIAS3_SIG, BIAS4_SIG, BIAS5_SIG, BIAS6_SIG, BIAS7_SIG, BIAS8_SIG, BIAS9_SIG : std_logic_vector(WIDTH+WIDTH-1 downto 0) := (others => '0');

begin

SET_O_VM <= SET_CNT;

DIN0_SIG   <= DIN0;
DIN1_SIG   <= DIN1;
DIN2_SIG   <= DIN2;
DIN3_SIG   <= DIN3;
DIN4_SIG   <= DIN4;
DIN5_SIG   <= DIN5;
DIN6_SIG   <= DIN6;
DIN7_SIG   <= DIN7;
DIN8_SIG   <= DIN8;
DIN9_SIG   <= DIN9;
DIN10_SIG  <= DIN10;
DIN11_SIG  <= DIN11;
DIN12_SIG  <= DIN12;
DIN13_SIG  <= DIN13;
DIN14_SIG  <= DIN14;
DIN15_SIG  <= DIN15;
DIN16_SIG  <= DIN16;
DIN17_SIG  <= DIN17;
DIN18_SIG  <= DIN18;
DIN19_SIG  <= DIN19;
DIN20_SIG  <= DIN20;
DIN21_SIG  <= DIN21;
DIN22_SIG  <= DIN22;
DIN23_SIG  <= DIN23;
DIN24_SIG  <= DIN24;
DIN25_SIG  <= DIN25;
DIN26_SIG  <= DIN26;
DIN27_SIG  <= DIN27;
DIN28_SIG  <= DIN28;
DIN29_SIG  <= DIN29;

O_VM0_INST: OUTPUT_VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER => 5)
Port map (
    CLK         =>  CLK,
    RESET       =>  RESET,
    SET         =>  SET_O_VM,
    DIN0        =>  DIN0_SIG,
    DIN1        =>  DIN1_SIG,
    DIN2        =>  DIN2_SIG,
    DIN3        =>  DIN3_SIG,
    DIN4        =>  DIN4_SIG,
    DIN5        =>  DIN5_SIG,
    DIN6        =>  DIN6_SIG,
    DIN7        =>  DIN7_SIG,
    DIN8        =>  DIN8_SIG,
    DIN9        =>  DIN9_SIG,
    DIN10       =>  DIN10_SIG,
    DIN11       =>  DIN11_SIG,
    DIN12       =>  DIN12_SIG,
    DIN13       =>  DIN13_SIG,
    DIN14       =>  DIN14_SIG,
    DIN15       =>  DIN15_SIG,
    DIN16       =>  DIN16_SIG,
    DIN17       =>  DIN17_SIG,
    DIN18       =>  DIN18_SIG,
    DIN19       =>  DIN19_SIG,
    DIN20       =>  DIN20_SIG,
    DIN21       =>  DIN21_SIG,
    DIN22       =>  DIN22_SIG,
    DIN23       =>  DIN23_SIG,
    DIN24       =>  DIN24_SIG,
    DIN25       =>  DIN25_SIG,
    DIN26       =>  DIN26_SIG,
    DIN27       =>  DIN27_SIG,
    DIN28       =>  DIN28_SIG,
    DIN29       =>  DIN29_SIG,
    ROM0_DATA   =>  ROM0_DATA0_SIG,
    ROM1_DATA   =>  ROM0_DATA1_SIG,
    ROM2_DATA   =>  ROM0_DATA2_SIG,
    ROM3_DATA   =>  ROM0_DATA3_SIG,
    ROM4_DATA   =>  ROM0_DATA4_SIG,
    ROM5_DATA   =>  ROM0_DATA5_SIG,
    ROM6_DATA   =>  ROM0_DATA6_SIG,
    ROM7_DATA   =>  ROM0_DATA7_SIG,
    ROM8_DATA   =>  ROM0_DATA8_SIG,
    ROM9_DATA   =>  ROM0_DATA9_SIG,
    ROM10_DATA  =>  ROM0_DATA10_SIG,
    ROM11_DATA  =>  ROM0_DATA11_SIG,
    ROM12_DATA  =>  ROM0_DATA12_SIG,
    ROM13_DATA  =>  ROM0_DATA13_SIG,
    ROM14_DATA  =>  ROM0_DATA14_SIG,
    ROM15_DATA  =>  ROM0_DATA15_SIG,
    ROM16_DATA  =>  ROM0_DATA16_SIG,
    ROM17_DATA  =>  ROM0_DATA17_SIG,
    ROM18_DATA  =>  ROM0_DATA18_SIG,
    ROM19_DATA  =>  ROM0_DATA19_SIG,
    ROM20_DATA  =>  ROM0_DATA20_SIG,
    ROM21_DATA  =>  ROM0_DATA21_SIG,
    ROM22_DATA  =>  ROM0_DATA22_SIG,
    ROM23_DATA  =>  ROM0_DATA23_SIG,
    ROM24_DATA  =>  ROM0_DATA24_SIG,
    ROM25_DATA  =>  ROM0_DATA25_SIG,
    ROM26_DATA  =>  ROM0_DATA26_SIG,
    ROM27_DATA  =>  ROM0_DATA27_SIG,
    ROM28_DATA  =>  ROM0_DATA28_SIG,
    ROM29_DATA  =>  ROM0_DATA29_SIG,
    ADDR0       =>  ADDR0_0_SIG,
    ADDR1       =>  ADDR0_1_SIG,
    ADDR2       =>  ADDR0_2_SIG,
    ADDR3       =>  ADDR0_3_SIG,
    ADDR4       =>  ADDR0_4_SIG,
    ADDR5       =>  ADDR0_5_SIG,
    ADDR6       =>  ADDR0_6_SIG,
    ADDR7       =>  ADDR0_7_SIG,
    ADDR8       =>  ADDR0_8_SIG,
    ADDR9       =>  ADDR0_9_SIG,
    ADDR10      =>  ADDR0_10_SIG,
    ADDR11      =>  ADDR0_11_SIG,
    ADDR12      =>  ADDR0_12_SIG,
    ADDR13      =>  ADDR0_13_SIG,
    ADDR14      =>  ADDR0_14_SIG,
    ADDR15      =>  ADDR0_15_SIG,
    ADDR16      =>  ADDR0_16_SIG,
    ADDR17      =>  ADDR0_17_SIG,
    ADDR18      =>  ADDR0_18_SIG,
    ADDR19      =>  ADDR0_19_SIG,
    ADDR20      =>  ADDR0_20_SIG,
    ADDR21      =>  ADDR0_21_SIG,
    ADDR22      =>  ADDR0_22_SIG,
    ADDR23      =>  ADDR0_23_SIG,
    ADDR24      =>  ADDR0_24_SIG,
    ADDR25      =>  ADDR0_25_SIG,
    ADDR26      =>  ADDR0_26_SIG,
    ADDR27      =>  ADDR0_27_SIG,
    ADDR28      =>  ADDR0_28_SIG,
    ADDR29      =>  ADDR0_29_SIG,
    DOUT        =>  O_VM0_OUT_SIG
);

O_VM1_INST: OUTPUT_VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER => 5)
Port map (
    CLK         =>  CLK,
    RESET       =>  RESET,
    SET         =>  SET_O_VM,
    DIN0        =>  DIN0_SIG,
    DIN1        =>  DIN1_SIG,
    DIN2        =>  DIN2_SIG,
    DIN3        =>  DIN3_SIG,
    DIN4        =>  DIN4_SIG,
    DIN5        =>  DIN5_SIG,
    DIN6        =>  DIN6_SIG,
    DIN7        =>  DIN7_SIG,
    DIN8        =>  DIN8_SIG,
    DIN9        =>  DIN9_SIG,
    DIN10       =>  DIN10_SIG,
    DIN11       =>  DIN11_SIG,
    DIN12       =>  DIN12_SIG,
    DIN13       =>  DIN13_SIG,
    DIN14       =>  DIN14_SIG,
    DIN15       =>  DIN15_SIG,
    DIN16       =>  DIN16_SIG,
    DIN17       =>  DIN17_SIG,
    DIN18       =>  DIN18_SIG,
    DIN19       =>  DIN19_SIG,
    DIN20       =>  DIN20_SIG,
    DIN21       =>  DIN21_SIG,
    DIN22       =>  DIN22_SIG,
    DIN23       =>  DIN23_SIG,
    DIN24       =>  DIN24_SIG,
    DIN25       =>  DIN25_SIG,
    DIN26       =>  DIN26_SIG,
    DIN27       =>  DIN27_SIG,
    DIN28       =>  DIN28_SIG,
    DIN29       =>  DIN29_SIG,
    ROM0_DATA   =>  ROM1_DATA0_SIG,
    ROM1_DATA   =>  ROM1_DATA1_SIG,
    ROM2_DATA   =>  ROM1_DATA2_SIG,
    ROM3_DATA   =>  ROM1_DATA3_SIG,
    ROM4_DATA   =>  ROM1_DATA4_SIG,
    ROM5_DATA   =>  ROM1_DATA5_SIG,
    ROM6_DATA   =>  ROM1_DATA6_SIG,
    ROM7_DATA   =>  ROM1_DATA7_SIG,
    ROM8_DATA   =>  ROM1_DATA8_SIG,
    ROM9_DATA   =>  ROM1_DATA9_SIG,
    ROM10_DATA  =>  ROM1_DATA10_SIG,
    ROM11_DATA  =>  ROM1_DATA11_SIG,
    ROM12_DATA  =>  ROM1_DATA12_SIG,
    ROM13_DATA  =>  ROM1_DATA13_SIG,
    ROM14_DATA  =>  ROM1_DATA14_SIG,
    ROM15_DATA  =>  ROM1_DATA15_SIG,
    ROM16_DATA  =>  ROM1_DATA16_SIG,
    ROM17_DATA  =>  ROM1_DATA17_SIG,
    ROM18_DATA  =>  ROM1_DATA18_SIG,
    ROM19_DATA  =>  ROM1_DATA19_SIG,
    ROM20_DATA  =>  ROM1_DATA20_SIG,
    ROM21_DATA  =>  ROM1_DATA21_SIG,
    ROM22_DATA  =>  ROM1_DATA22_SIG,
    ROM23_DATA  =>  ROM1_DATA23_SIG,
    ROM24_DATA  =>  ROM1_DATA24_SIG,
    ROM25_DATA  =>  ROM1_DATA25_SIG,
    ROM26_DATA  =>  ROM1_DATA26_SIG,
    ROM27_DATA  =>  ROM1_DATA27_SIG,
    ROM28_DATA  =>  ROM1_DATA28_SIG,
    ROM29_DATA  =>  ROM0_DATA29_SIG,
    ADDR0       =>  ADDR1_0_SIG,
    ADDR1       =>  ADDR1_1_SIG,
    ADDR2       =>  ADDR1_2_SIG,
    ADDR3       =>  ADDR1_3_SIG,
    ADDR4       =>  ADDR1_4_SIG,
    ADDR5       =>  ADDR1_5_SIG,
    ADDR6       =>  ADDR1_6_SIG,
    ADDR7       =>  ADDR1_7_SIG,
    ADDR8       =>  ADDR1_8_SIG,
    ADDR9       =>  ADDR1_9_SIG,
    ADDR10      =>  ADDR1_10_SIG,
    ADDR11      =>  ADDR1_11_SIG,
    ADDR12      =>  ADDR1_12_SIG,
    ADDR13      =>  ADDR1_13_SIG,
    ADDR14      =>  ADDR1_14_SIG,
    ADDR15      =>  ADDR1_15_SIG,
    ADDR16      =>  ADDR1_16_SIG,
    ADDR17      =>  ADDR1_17_SIG,
    ADDR18      =>  ADDR1_18_SIG,
    ADDR19      =>  ADDR1_19_SIG,
    ADDR20      =>  ADDR1_20_SIG,
    ADDR21      =>  ADDR1_21_SIG,
    ADDR22      =>  ADDR1_22_SIG,
    ADDR23      =>  ADDR1_23_SIG,
    ADDR24      =>  ADDR1_24_SIG,
    ADDR25      =>  ADDR1_25_SIG,
    ADDR26      =>  ADDR1_26_SIG,
    ADDR27      =>  ADDR1_27_SIG,
    ADDR28      =>  ADDR1_28_SIG,
    ADDR29      =>  ADDR1_29_SIG,
    DOUT        =>  O_VM1_OUT_SIG
);

O_VM2_INST: OUTPUT_VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER => 5)
Port map (
    CLK         =>  CLK,
    RESET       =>  RESET,
    SET         =>  SET_O_VM,
    DIN0        =>  DIN0_SIG,
    DIN1        =>  DIN1_SIG,
    DIN2        =>  DIN2_SIG,
    DIN3        =>  DIN3_SIG,
    DIN4        =>  DIN4_SIG,
    DIN5        =>  DIN5_SIG,
    DIN6        =>  DIN6_SIG,
    DIN7        =>  DIN7_SIG,
    DIN8        =>  DIN8_SIG,
    DIN9        =>  DIN9_SIG,
    DIN10       =>  DIN10_SIG,
    DIN11       =>  DIN11_SIG,
    DIN12       =>  DIN12_SIG,
    DIN13       =>  DIN13_SIG,
    DIN14       =>  DIN14_SIG,
    DIN15       =>  DIN15_SIG,
    DIN16       =>  DIN16_SIG,
    DIN17       =>  DIN17_SIG,
    DIN18       =>  DIN18_SIG,
    DIN19       =>  DIN19_SIG,
    DIN20       =>  DIN20_SIG,
    DIN21       =>  DIN21_SIG,
    DIN22       =>  DIN22_SIG,
    DIN23       =>  DIN23_SIG,
    DIN24       =>  DIN24_SIG,
    DIN25       =>  DIN25_SIG,
    DIN26       =>  DIN26_SIG,
    DIN27       =>  DIN27_SIG,
    DIN28       =>  DIN28_SIG,
    DIN29       =>  DIN29_SIG,
    ROM0_DATA   =>  ROM2_DATA0_SIG,
    ROM1_DATA   =>  ROM2_DATA1_SIG,
    ROM2_DATA   =>  ROM2_DATA2_SIG,
    ROM3_DATA   =>  ROM2_DATA3_SIG,
    ROM4_DATA   =>  ROM2_DATA4_SIG,
    ROM5_DATA   =>  ROM2_DATA5_SIG,
    ROM6_DATA   =>  ROM2_DATA6_SIG,
    ROM7_DATA   =>  ROM2_DATA7_SIG,
    ROM8_DATA   =>  ROM2_DATA8_SIG,
    ROM9_DATA   =>  ROM2_DATA9_SIG,
    ROM10_DATA  =>  ROM2_DATA10_SIG,
    ROM11_DATA  =>  ROM2_DATA11_SIG,
    ROM12_DATA  =>  ROM2_DATA12_SIG,
    ROM13_DATA  =>  ROM2_DATA13_SIG,
    ROM14_DATA  =>  ROM2_DATA14_SIG,
    ROM15_DATA  =>  ROM2_DATA15_SIG,
    ROM16_DATA  =>  ROM2_DATA16_SIG,
    ROM17_DATA  =>  ROM2_DATA17_SIG,
    ROM18_DATA  =>  ROM2_DATA18_SIG,
    ROM19_DATA  =>  ROM2_DATA19_SIG,
    ROM20_DATA  =>  ROM2_DATA20_SIG,
    ROM21_DATA  =>  ROM2_DATA21_SIG,
    ROM22_DATA  =>  ROM2_DATA22_SIG,
    ROM23_DATA  =>  ROM2_DATA23_SIG,
    ROM24_DATA  =>  ROM2_DATA24_SIG,
    ROM25_DATA  =>  ROM2_DATA25_SIG,
    ROM26_DATA  =>  ROM2_DATA26_SIG,
    ROM27_DATA  =>  ROM2_DATA27_SIG,
    ROM28_DATA  =>  ROM2_DATA28_SIG,
    ROM29_DATA  =>  ROM2_DATA29_SIG,
    ADDR0       =>  ADDR2_0_SIG,
    ADDR1       =>  ADDR2_1_SIG,
    ADDR2       =>  ADDR2_2_SIG,
    ADDR3       =>  ADDR2_3_SIG,
    ADDR4       =>  ADDR2_4_SIG,
    ADDR5       =>  ADDR2_5_SIG,
    ADDR6       =>  ADDR2_6_SIG,
    ADDR7       =>  ADDR2_7_SIG,
    ADDR8       =>  ADDR2_8_SIG,
    ADDR9       =>  ADDR2_9_SIG,
    ADDR10      =>  ADDR2_10_SIG,
    ADDR11      =>  ADDR2_11_SIG,
    ADDR12      =>  ADDR2_12_SIG,
    ADDR13      =>  ADDR2_13_SIG,
    ADDR14      =>  ADDR2_14_SIG,
    ADDR15      =>  ADDR2_15_SIG,
    ADDR16      =>  ADDR2_16_SIG,
    ADDR17      =>  ADDR2_17_SIG,
    ADDR18      =>  ADDR2_18_SIG,
    ADDR19      =>  ADDR2_19_SIG,
    ADDR20      =>  ADDR2_20_SIG,
    ADDR21      =>  ADDR2_21_SIG,
    ADDR22      =>  ADDR2_22_SIG,
    ADDR23      =>  ADDR2_23_SIG,
    ADDR24      =>  ADDR2_24_SIG,
    ADDR25      =>  ADDR2_25_SIG,
    ADDR26      =>  ADDR2_26_SIG,
    ADDR27      =>  ADDR2_27_SIG,
    ADDR28      =>  ADDR2_28_SIG,
    ADDR29      =>  ADDR2_29_SIG,
    DOUT        =>  O_VM2_OUT_SIG
);

O_VM3_INST: OUTPUT_VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER => 5)
Port map (
    CLK         =>  CLK,
    RESET       =>  RESET,
    SET         =>  SET_O_VM,
    DIN0        =>  DIN0_SIG,
    DIN1        =>  DIN1_SIG,
    DIN2        =>  DIN2_SIG,
    DIN3        =>  DIN3_SIG,
    DIN4        =>  DIN4_SIG,
    DIN5        =>  DIN5_SIG,
    DIN6        =>  DIN6_SIG,
    DIN7        =>  DIN7_SIG,
    DIN8        =>  DIN8_SIG,
    DIN9        =>  DIN9_SIG,
    DIN10       =>  DIN10_SIG,
    DIN11       =>  DIN11_SIG,
    DIN12       =>  DIN12_SIG,
    DIN13       =>  DIN13_SIG,
    DIN14       =>  DIN14_SIG,
    DIN15       =>  DIN15_SIG,
    DIN16       =>  DIN16_SIG,
    DIN17       =>  DIN17_SIG,
    DIN18       =>  DIN18_SIG,
    DIN19       =>  DIN19_SIG,
    DIN20       =>  DIN20_SIG,
    DIN21       =>  DIN21_SIG,
    DIN22       =>  DIN22_SIG,
    DIN23       =>  DIN23_SIG,
    DIN24       =>  DIN24_SIG,
    DIN25       =>  DIN25_SIG,
    DIN26       =>  DIN26_SIG,
    DIN27       =>  DIN27_SIG,
    DIN28       =>  DIN28_SIG,
    DIN29       =>  DIN29_SIG,
    ROM0_DATA   =>  ROM3_DATA0_SIG,
    ROM1_DATA   =>  ROM3_DATA1_SIG,
    ROM2_DATA   =>  ROM3_DATA2_SIG,
    ROM3_DATA   =>  ROM3_DATA3_SIG,
    ROM4_DATA   =>  ROM3_DATA4_SIG,
    ROM5_DATA   =>  ROM3_DATA5_SIG,
    ROM6_DATA   =>  ROM3_DATA6_SIG,
    ROM7_DATA   =>  ROM3_DATA7_SIG,
    ROM8_DATA   =>  ROM3_DATA8_SIG,
    ROM9_DATA   =>  ROM3_DATA9_SIG,
    ROM10_DATA  =>  ROM3_DATA10_SIG,
    ROM11_DATA  =>  ROM3_DATA11_SIG,
    ROM12_DATA  =>  ROM3_DATA12_SIG,
    ROM13_DATA  =>  ROM3_DATA13_SIG,
    ROM14_DATA  =>  ROM3_DATA14_SIG,
    ROM15_DATA  =>  ROM3_DATA15_SIG,
    ROM16_DATA  =>  ROM3_DATA16_SIG,
    ROM17_DATA  =>  ROM3_DATA17_SIG,
    ROM18_DATA  =>  ROM3_DATA18_SIG,
    ROM19_DATA  =>  ROM3_DATA19_SIG,
    ROM20_DATA  =>  ROM3_DATA20_SIG,
    ROM21_DATA  =>  ROM3_DATA21_SIG,
    ROM22_DATA  =>  ROM3_DATA22_SIG,
    ROM23_DATA  =>  ROM3_DATA23_SIG,
    ROM24_DATA  =>  ROM3_DATA24_SIG,
    ROM25_DATA  =>  ROM3_DATA25_SIG,
    ROM26_DATA  =>  ROM3_DATA26_SIG,
    ROM27_DATA  =>  ROM3_DATA27_SIG,
    ROM28_DATA  =>  ROM3_DATA28_SIG,
    ROM29_DATA  =>  ROM3_DATA29_SIG,
    ADDR0       =>  ADDR3_0_SIG,
    ADDR1       =>  ADDR3_1_SIG,
    ADDR2       =>  ADDR3_2_SIG,
    ADDR3       =>  ADDR3_3_SIG,
    ADDR4       =>  ADDR3_4_SIG,
    ADDR5       =>  ADDR3_5_SIG,
    ADDR6       =>  ADDR3_6_SIG,
    ADDR7       =>  ADDR3_7_SIG,
    ADDR8       =>  ADDR3_8_SIG,
    ADDR9       =>  ADDR3_9_SIG,
    ADDR10      =>  ADDR3_10_SIG,
    ADDR11      =>  ADDR3_11_SIG,
    ADDR12      =>  ADDR3_12_SIG,
    ADDR13      =>  ADDR3_13_SIG,
    ADDR14      =>  ADDR3_14_SIG,
    ADDR15      =>  ADDR3_15_SIG,
    ADDR16      =>  ADDR3_16_SIG,
    ADDR17      =>  ADDR3_17_SIG,
    ADDR18      =>  ADDR3_18_SIG,
    ADDR19      =>  ADDR3_19_SIG,
    ADDR20      =>  ADDR3_20_SIG,
    ADDR21      =>  ADDR3_21_SIG,
    ADDR22      =>  ADDR3_22_SIG,
    ADDR23      =>  ADDR3_23_SIG,
    ADDR24      =>  ADDR3_24_SIG,
    ADDR25      =>  ADDR3_25_SIG,
    ADDR26      =>  ADDR3_26_SIG,
    ADDR27      =>  ADDR3_27_SIG,
    ADDR28      =>  ADDR3_28_SIG,
    ADDR29      =>  ADDR3_29_SIG,
    DOUT        =>  O_VM3_OUT_SIG
);

O_VM4_INST: OUTPUT_VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER => 5)
Port map (
    CLK         =>  CLK,
    RESET       =>  RESET,
    SET         =>  SET_O_VM,
    DIN0        =>  DIN0_SIG,
    DIN1        =>  DIN1_SIG,
    DIN2        =>  DIN2_SIG,
    DIN3        =>  DIN3_SIG,
    DIN4        =>  DIN4_SIG,
    DIN5        =>  DIN5_SIG,
    DIN6        =>  DIN6_SIG,
    DIN7        =>  DIN7_SIG,
    DIN8        =>  DIN8_SIG,
    DIN9        =>  DIN9_SIG,
    DIN10       =>  DIN10_SIG,
    DIN11       =>  DIN11_SIG,
    DIN12       =>  DIN12_SIG,
    DIN13       =>  DIN13_SIG,
    DIN14       =>  DIN14_SIG,
    DIN15       =>  DIN15_SIG,
    DIN16       =>  DIN16_SIG,
    DIN17       =>  DIN17_SIG,
    DIN18       =>  DIN18_SIG,
    DIN19       =>  DIN19_SIG,
    DIN20       =>  DIN20_SIG,
    DIN21       =>  DIN21_SIG,
    DIN22       =>  DIN22_SIG,
    DIN23       =>  DIN23_SIG,
    DIN24       =>  DIN24_SIG,
    DIN25       =>  DIN25_SIG,
    DIN26       =>  DIN26_SIG,
    DIN27       =>  DIN27_SIG,
    DIN28       =>  DIN28_SIG,
    DIN29       =>  DIN29_SIG,
    ROM0_DATA   =>  ROM4_DATA0_SIG,
    ROM1_DATA   =>  ROM4_DATA1_SIG,
    ROM2_DATA   =>  ROM4_DATA2_SIG,
    ROM3_DATA   =>  ROM4_DATA3_SIG,
    ROM4_DATA   =>  ROM4_DATA4_SIG,
    ROM5_DATA   =>  ROM4_DATA5_SIG,
    ROM6_DATA   =>  ROM4_DATA6_SIG,
    ROM7_DATA   =>  ROM4_DATA7_SIG,
    ROM8_DATA   =>  ROM4_DATA8_SIG,
    ROM9_DATA   =>  ROM4_DATA9_SIG,
    ROM10_DATA  =>  ROM4_DATA10_SIG,
    ROM11_DATA  =>  ROM4_DATA11_SIG,
    ROM12_DATA  =>  ROM4_DATA12_SIG,
    ROM13_DATA  =>  ROM4_DATA13_SIG,
    ROM14_DATA  =>  ROM4_DATA14_SIG,
    ROM15_DATA  =>  ROM4_DATA15_SIG,
    ROM16_DATA  =>  ROM4_DATA16_SIG,
    ROM17_DATA  =>  ROM4_DATA17_SIG,
    ROM18_DATA  =>  ROM4_DATA18_SIG,
    ROM19_DATA  =>  ROM4_DATA19_SIG,
    ROM20_DATA  =>  ROM4_DATA20_SIG,
    ROM21_DATA  =>  ROM4_DATA21_SIG,
    ROM22_DATA  =>  ROM4_DATA22_SIG,
    ROM23_DATA  =>  ROM4_DATA23_SIG,
    ROM24_DATA  =>  ROM4_DATA24_SIG,
    ROM25_DATA  =>  ROM4_DATA25_SIG,
    ROM26_DATA  =>  ROM4_DATA26_SIG,
    ROM27_DATA  =>  ROM4_DATA27_SIG,
    ROM28_DATA  =>  ROM4_DATA28_SIG,
    ROM29_DATA  =>  ROM4_DATA29_SIG,
    ADDR0       =>  ADDR4_0_SIG,
    ADDR1       =>  ADDR4_1_SIG,
    ADDR2       =>  ADDR4_2_SIG,
    ADDR3       =>  ADDR4_3_SIG,
    ADDR4       =>  ADDR4_4_SIG,
    ADDR5       =>  ADDR4_5_SIG,
    ADDR6       =>  ADDR4_6_SIG,
    ADDR7       =>  ADDR4_7_SIG,
    ADDR8       =>  ADDR4_8_SIG,
    ADDR9       =>  ADDR4_9_SIG,
    ADDR10      =>  ADDR4_10_SIG,
    ADDR11      =>  ADDR4_11_SIG,
    ADDR12      =>  ADDR4_12_SIG,
    ADDR13      =>  ADDR4_13_SIG,
    ADDR14      =>  ADDR4_14_SIG,
    ADDR15      =>  ADDR4_15_SIG,
    ADDR16      =>  ADDR4_16_SIG,
    ADDR17      =>  ADDR4_17_SIG,
    ADDR18      =>  ADDR4_18_SIG,
    ADDR19      =>  ADDR4_19_SIG,
    ADDR20      =>  ADDR4_20_SIG,
    ADDR21      =>  ADDR4_21_SIG,
    ADDR22      =>  ADDR4_22_SIG,
    ADDR23      =>  ADDR4_23_SIG,
    ADDR24      =>  ADDR4_24_SIG,
    ADDR25      =>  ADDR4_25_SIG,
    ADDR26      =>  ADDR4_26_SIG,
    ADDR27      =>  ADDR4_27_SIG,
    ADDR28      =>  ADDR4_28_SIG,
    ADDR29      =>  ADDR4_29_SIG,
    DOUT        =>  O_VM4_OUT_SIG
);

O_VM5_INST: OUTPUT_VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER => 5)
Port map (
    CLK         =>  CLK,
    RESET       =>  RESET,
    SET         =>  SET_O_VM,
    DIN0        =>  DIN0_SIG,
    DIN1        =>  DIN1_SIG,
    DIN2        =>  DIN2_SIG,
    DIN3        =>  DIN3_SIG,
    DIN4        =>  DIN4_SIG,
    DIN5        =>  DIN5_SIG,
    DIN6        =>  DIN6_SIG,
    DIN7        =>  DIN7_SIG,
    DIN8        =>  DIN8_SIG,
    DIN9        =>  DIN9_SIG,
    DIN10       =>  DIN10_SIG,
    DIN11       =>  DIN11_SIG,
    DIN12       =>  DIN12_SIG,
    DIN13       =>  DIN13_SIG,
    DIN14       =>  DIN14_SIG,
    DIN15       =>  DIN15_SIG,
    DIN16       =>  DIN16_SIG,
    DIN17       =>  DIN17_SIG,
    DIN18       =>  DIN18_SIG,
    DIN19       =>  DIN19_SIG,
    DIN20       =>  DIN20_SIG,
    DIN21       =>  DIN21_SIG,
    DIN22       =>  DIN22_SIG,
    DIN23       =>  DIN23_SIG,
    DIN24       =>  DIN24_SIG,
    DIN25       =>  DIN25_SIG,
    DIN26       =>  DIN26_SIG,
    DIN27       =>  DIN27_SIG,
    DIN28       =>  DIN28_SIG,
    DIN29       =>  DIN29_SIG,
    ROM0_DATA   =>  ROM5_DATA0_SIG,
    ROM1_DATA   =>  ROM5_DATA1_SIG,
    ROM2_DATA   =>  ROM5_DATA2_SIG,
    ROM3_DATA   =>  ROM5_DATA3_SIG,
    ROM4_DATA   =>  ROM5_DATA4_SIG,
    ROM5_DATA   =>  ROM5_DATA5_SIG,
    ROM6_DATA   =>  ROM5_DATA6_SIG,
    ROM7_DATA   =>  ROM5_DATA7_SIG,
    ROM8_DATA   =>  ROM5_DATA8_SIG,
    ROM9_DATA   =>  ROM5_DATA9_SIG,
    ROM10_DATA  =>  ROM5_DATA10_SIG,
    ROM11_DATA  =>  ROM5_DATA11_SIG,
    ROM12_DATA  =>  ROM5_DATA12_SIG,
    ROM13_DATA  =>  ROM5_DATA13_SIG,
    ROM14_DATA  =>  ROM5_DATA14_SIG,
    ROM15_DATA  =>  ROM5_DATA15_SIG,
    ROM16_DATA  =>  ROM5_DATA16_SIG,
    ROM17_DATA  =>  ROM5_DATA17_SIG,
    ROM18_DATA  =>  ROM5_DATA18_SIG,
    ROM19_DATA  =>  ROM5_DATA19_SIG,
    ROM20_DATA  =>  ROM5_DATA20_SIG,
    ROM21_DATA  =>  ROM5_DATA21_SIG,
    ROM22_DATA  =>  ROM5_DATA22_SIG,
    ROM23_DATA  =>  ROM5_DATA23_SIG,
    ROM24_DATA  =>  ROM5_DATA24_SIG,
    ROM25_DATA  =>  ROM5_DATA25_SIG,
    ROM26_DATA  =>  ROM5_DATA26_SIG,
    ROM27_DATA  =>  ROM5_DATA27_SIG,
    ROM28_DATA  =>  ROM5_DATA28_SIG,
    ROM29_DATA  =>  ROM5_DATA29_SIG,
    ADDR0       =>  ADDR5_0_SIG,
    ADDR1       =>  ADDR5_1_SIG,
    ADDR2       =>  ADDR5_2_SIG,
    ADDR3       =>  ADDR5_3_SIG,
    ADDR4       =>  ADDR5_4_SIG,
    ADDR5       =>  ADDR5_5_SIG,
    ADDR6       =>  ADDR5_6_SIG,
    ADDR7       =>  ADDR5_7_SIG,
    ADDR8       =>  ADDR5_8_SIG,
    ADDR9       =>  ADDR5_9_SIG,
    ADDR10      =>  ADDR5_10_SIG,
    ADDR11      =>  ADDR5_11_SIG,
    ADDR12      =>  ADDR5_12_SIG,
    ADDR13      =>  ADDR5_13_SIG,
    ADDR14      =>  ADDR5_14_SIG,
    ADDR15      =>  ADDR5_15_SIG,
    ADDR16      =>  ADDR5_16_SIG,
    ADDR17      =>  ADDR5_17_SIG,
    ADDR18      =>  ADDR5_18_SIG,
    ADDR19      =>  ADDR5_19_SIG,
    ADDR20      =>  ADDR5_20_SIG,
    ADDR21      =>  ADDR5_21_SIG,
    ADDR22      =>  ADDR5_22_SIG,
    ADDR23      =>  ADDR5_23_SIG,
    ADDR24      =>  ADDR5_24_SIG,
    ADDR25      =>  ADDR5_25_SIG,
    ADDR26      =>  ADDR5_26_SIG,
    ADDR27      =>  ADDR5_27_SIG,
    ADDR28      =>  ADDR5_28_SIG,
    ADDR29      =>  ADDR5_29_SIG,
    DOUT        =>  O_VM5_OUT_SIG
);

O_VM6_INST: OUTPUT_VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER => 5)
Port map (
    CLK         =>  CLK,
    RESET       =>  RESET,
    SET         =>  SET_O_VM,
    DIN0        =>  DIN0_SIG,
    DIN1        =>  DIN1_SIG,
    DIN2        =>  DIN2_SIG,
    DIN3        =>  DIN3_SIG,
    DIN4        =>  DIN4_SIG,
    DIN5        =>  DIN5_SIG,
    DIN6        =>  DIN6_SIG,
    DIN7        =>  DIN7_SIG,
    DIN8        =>  DIN8_SIG,
    DIN9        =>  DIN9_SIG,
    DIN10       =>  DIN10_SIG,
    DIN11       =>  DIN11_SIG,
    DIN12       =>  DIN12_SIG,
    DIN13       =>  DIN13_SIG,
    DIN14       =>  DIN14_SIG,
    DIN15       =>  DIN15_SIG,
    DIN16       =>  DIN16_SIG,
    DIN17       =>  DIN17_SIG,
    DIN18       =>  DIN18_SIG,
    DIN19       =>  DIN19_SIG,
    DIN20       =>  DIN20_SIG,
    DIN21       =>  DIN21_SIG,
    DIN22       =>  DIN22_SIG,
    DIN23       =>  DIN23_SIG,
    DIN24       =>  DIN24_SIG,
    DIN25       =>  DIN25_SIG,
    DIN26       =>  DIN26_SIG,
    DIN27       =>  DIN27_SIG,
    DIN28       =>  DIN28_SIG,
    DIN29       =>  DIN29_SIG,
    ROM0_DATA   =>  ROM6_DATA0_SIG,
    ROM1_DATA   =>  ROM6_DATA1_SIG,
    ROM2_DATA   =>  ROM6_DATA2_SIG,
    ROM3_DATA   =>  ROM6_DATA3_SIG,
    ROM4_DATA   =>  ROM6_DATA4_SIG,
    ROM5_DATA   =>  ROM6_DATA5_SIG,
    ROM6_DATA   =>  ROM6_DATA6_SIG,
    ROM7_DATA   =>  ROM6_DATA7_SIG,
    ROM8_DATA   =>  ROM6_DATA8_SIG,
    ROM9_DATA   =>  ROM6_DATA9_SIG,
    ROM10_DATA  =>  ROM6_DATA10_SIG,
    ROM11_DATA  =>  ROM6_DATA11_SIG,
    ROM12_DATA  =>  ROM6_DATA12_SIG,
    ROM13_DATA  =>  ROM6_DATA13_SIG,
    ROM14_DATA  =>  ROM6_DATA14_SIG,
    ROM15_DATA  =>  ROM6_DATA15_SIG,
    ROM16_DATA  =>  ROM6_DATA16_SIG,
    ROM17_DATA  =>  ROM6_DATA17_SIG,
    ROM18_DATA  =>  ROM6_DATA18_SIG,
    ROM19_DATA  =>  ROM6_DATA19_SIG,
    ROM20_DATA  =>  ROM6_DATA20_SIG,
    ROM21_DATA  =>  ROM6_DATA21_SIG,
    ROM22_DATA  =>  ROM6_DATA22_SIG,
    ROM23_DATA  =>  ROM6_DATA23_SIG,
    ROM24_DATA  =>  ROM6_DATA24_SIG,
    ROM25_DATA  =>  ROM6_DATA25_SIG,
    ROM26_DATA  =>  ROM6_DATA26_SIG,
    ROM27_DATA  =>  ROM6_DATA27_SIG,
    ROM28_DATA  =>  ROM6_DATA28_SIG,
    ROM29_DATA  =>  ROM6_DATA29_SIG,
    ADDR0       =>  ADDR6_0_SIG,
    ADDR1       =>  ADDR6_1_SIG,
    ADDR2       =>  ADDR6_2_SIG,
    ADDR3       =>  ADDR6_3_SIG,
    ADDR4       =>  ADDR6_4_SIG,
    ADDR5       =>  ADDR6_5_SIG,
    ADDR6       =>  ADDR6_6_SIG,
    ADDR7       =>  ADDR6_7_SIG,
    ADDR8       =>  ADDR6_8_SIG,
    ADDR9       =>  ADDR6_9_SIG,
    ADDR10      =>  ADDR6_10_SIG,
    ADDR11      =>  ADDR6_11_SIG,
    ADDR12      =>  ADDR6_12_SIG,
    ADDR13      =>  ADDR6_13_SIG,
    ADDR14      =>  ADDR6_14_SIG,
    ADDR15      =>  ADDR6_15_SIG,
    ADDR16      =>  ADDR6_16_SIG,
    ADDR17      =>  ADDR6_17_SIG,
    ADDR18      =>  ADDR6_18_SIG,
    ADDR19      =>  ADDR6_19_SIG,
    ADDR20      =>  ADDR6_20_SIG,
    ADDR21      =>  ADDR6_21_SIG,
    ADDR22      =>  ADDR6_22_SIG,
    ADDR23      =>  ADDR6_23_SIG,
    ADDR24      =>  ADDR6_24_SIG,
    ADDR25      =>  ADDR6_25_SIG,
    ADDR26      =>  ADDR6_26_SIG,
    ADDR27      =>  ADDR6_27_SIG,
    ADDR28      =>  ADDR6_28_SIG,
    ADDR29      =>  ADDR6_29_SIG,
    DOUT        =>  O_VM6_OUT_SIG
);

O_VM7_INST: OUTPUT_VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER => 5)
Port map (
    CLK         =>  CLK,
    RESET       =>  RESET,
    SET         =>  SET_O_VM,
    DIN0        =>  DIN0_SIG,
    DIN1        =>  DIN1_SIG,
    DIN2        =>  DIN2_SIG,
    DIN3        =>  DIN3_SIG,
    DIN4        =>  DIN4_SIG,
    DIN5        =>  DIN5_SIG,
    DIN6        =>  DIN6_SIG,
    DIN7        =>  DIN7_SIG,
    DIN8        =>  DIN8_SIG,
    DIN9        =>  DIN9_SIG,
    DIN10       =>  DIN10_SIG,
    DIN11       =>  DIN11_SIG,
    DIN12       =>  DIN12_SIG,
    DIN13       =>  DIN13_SIG,
    DIN14       =>  DIN14_SIG,
    DIN15       =>  DIN15_SIG,
    DIN16       =>  DIN16_SIG,
    DIN17       =>  DIN17_SIG,
    DIN18       =>  DIN18_SIG,
    DIN19       =>  DIN19_SIG,
    DIN20       =>  DIN20_SIG,
    DIN21       =>  DIN21_SIG,
    DIN22       =>  DIN22_SIG,
    DIN23       =>  DIN23_SIG,
    DIN24       =>  DIN24_SIG,
    DIN25       =>  DIN25_SIG,
    DIN26       =>  DIN26_SIG,
    DIN27       =>  DIN27_SIG,
    DIN28       =>  DIN28_SIG,
    DIN29       =>  DIN29_SIG,
    ROM0_DATA   =>  ROM7_DATA0_SIG,
    ROM1_DATA   =>  ROM7_DATA1_SIG,
    ROM2_DATA   =>  ROM7_DATA2_SIG,
    ROM3_DATA   =>  ROM7_DATA3_SIG,
    ROM4_DATA   =>  ROM7_DATA4_SIG,
    ROM5_DATA   =>  ROM7_DATA5_SIG,
    ROM6_DATA   =>  ROM7_DATA6_SIG,
    ROM7_DATA   =>  ROM7_DATA7_SIG,
    ROM8_DATA   =>  ROM7_DATA8_SIG,
    ROM9_DATA   =>  ROM7_DATA9_SIG,
    ROM10_DATA  =>  ROM7_DATA10_SIG,
    ROM11_DATA  =>  ROM7_DATA11_SIG,
    ROM12_DATA  =>  ROM7_DATA12_SIG,
    ROM13_DATA  =>  ROM7_DATA13_SIG,
    ROM14_DATA  =>  ROM7_DATA14_SIG,
    ROM15_DATA  =>  ROM7_DATA15_SIG,
    ROM16_DATA  =>  ROM7_DATA16_SIG,
    ROM17_DATA  =>  ROM7_DATA17_SIG,
    ROM18_DATA  =>  ROM7_DATA18_SIG,
    ROM19_DATA  =>  ROM7_DATA19_SIG,
    ROM20_DATA  =>  ROM7_DATA20_SIG,
    ROM21_DATA  =>  ROM7_DATA21_SIG,
    ROM22_DATA  =>  ROM7_DATA22_SIG,
    ROM23_DATA  =>  ROM7_DATA23_SIG,
    ROM24_DATA  =>  ROM7_DATA24_SIG,
    ROM25_DATA  =>  ROM7_DATA25_SIG,
    ROM26_DATA  =>  ROM7_DATA26_SIG,
    ROM27_DATA  =>  ROM7_DATA27_SIG,
    ROM28_DATA  =>  ROM7_DATA28_SIG,
    ROM29_DATA  =>  ROM7_DATA29_SIG,
    ADDR0       =>  ADDR7_0_SIG,
    ADDR1       =>  ADDR7_1_SIG,
    ADDR2       =>  ADDR7_2_SIG,
    ADDR3       =>  ADDR7_3_SIG,
    ADDR4       =>  ADDR7_4_SIG,
    ADDR5       =>  ADDR7_5_SIG,
    ADDR6       =>  ADDR7_6_SIG,
    ADDR7       =>  ADDR7_7_SIG,
    ADDR8       =>  ADDR7_8_SIG,
    ADDR9       =>  ADDR7_9_SIG,
    ADDR10      =>  ADDR7_10_SIG,
    ADDR11      =>  ADDR7_11_SIG,
    ADDR12      =>  ADDR7_12_SIG,
    ADDR13      =>  ADDR7_13_SIG,
    ADDR14      =>  ADDR7_14_SIG,
    ADDR15      =>  ADDR7_15_SIG,
    ADDR16      =>  ADDR7_16_SIG,
    ADDR17      =>  ADDR7_17_SIG,
    ADDR18      =>  ADDR7_18_SIG,
    ADDR19      =>  ADDR7_19_SIG,
    ADDR20      =>  ADDR7_20_SIG,
    ADDR21      =>  ADDR7_21_SIG,
    ADDR22      =>  ADDR7_22_SIG,
    ADDR23      =>  ADDR7_23_SIG,
    ADDR24      =>  ADDR7_24_SIG,
    ADDR25      =>  ADDR7_25_SIG,
    ADDR26      =>  ADDR7_26_SIG,
    ADDR27      =>  ADDR7_27_SIG,
    ADDR28      =>  ADDR7_28_SIG,
    ADDR29      =>  ADDR7_29_SIG,
    DOUT        =>  O_VM7_OUT_SIG
);

O_VM8_INST: OUTPUT_VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER => 5)
Port map (
    CLK         =>  CLK,
    RESET       =>  RESET,
    SET         =>  SET_O_VM,
    DIN0        =>  DIN0_SIG,
    DIN1        =>  DIN1_SIG,
    DIN2        =>  DIN2_SIG,
    DIN3        =>  DIN3_SIG,
    DIN4        =>  DIN4_SIG,
    DIN5        =>  DIN5_SIG,
    DIN6        =>  DIN6_SIG,
    DIN7        =>  DIN7_SIG,
    DIN8        =>  DIN8_SIG,
    DIN9        =>  DIN9_SIG,
    DIN10       =>  DIN10_SIG,
    DIN11       =>  DIN11_SIG,
    DIN12       =>  DIN12_SIG,
    DIN13       =>  DIN13_SIG,
    DIN14       =>  DIN14_SIG,
    DIN15       =>  DIN15_SIG,
    DIN16       =>  DIN16_SIG,
    DIN17       =>  DIN17_SIG,
    DIN18       =>  DIN18_SIG,
    DIN19       =>  DIN19_SIG,
    DIN20       =>  DIN20_SIG,
    DIN21       =>  DIN21_SIG,
    DIN22       =>  DIN22_SIG,
    DIN23       =>  DIN23_SIG,
    DIN24       =>  DIN24_SIG,
    DIN25       =>  DIN25_SIG,
    DIN26       =>  DIN26_SIG,
    DIN27       =>  DIN27_SIG,
    DIN28       =>  DIN28_SIG,
    DIN29       =>  DIN29_SIG,
    ROM0_DATA   =>  ROM8_DATA0_SIG,
    ROM1_DATA   =>  ROM8_DATA1_SIG,
    ROM2_DATA   =>  ROM8_DATA2_SIG,
    ROM3_DATA   =>  ROM8_DATA3_SIG,
    ROM4_DATA   =>  ROM8_DATA4_SIG,
    ROM5_DATA   =>  ROM8_DATA5_SIG,
    ROM6_DATA   =>  ROM8_DATA6_SIG,
    ROM7_DATA   =>  ROM8_DATA7_SIG,
    ROM8_DATA   =>  ROM8_DATA8_SIG,
    ROM9_DATA   =>  ROM8_DATA9_SIG,
    ROM10_DATA  =>  ROM8_DATA10_SIG,
    ROM11_DATA  =>  ROM8_DATA11_SIG,
    ROM12_DATA  =>  ROM8_DATA12_SIG,
    ROM13_DATA  =>  ROM8_DATA13_SIG,
    ROM14_DATA  =>  ROM8_DATA14_SIG,
    ROM15_DATA  =>  ROM8_DATA15_SIG,
    ROM16_DATA  =>  ROM8_DATA16_SIG,
    ROM17_DATA  =>  ROM8_DATA17_SIG,
    ROM18_DATA  =>  ROM8_DATA18_SIG,
    ROM19_DATA  =>  ROM8_DATA19_SIG,
    ROM20_DATA  =>  ROM8_DATA20_SIG,
    ROM21_DATA  =>  ROM8_DATA21_SIG,
    ROM22_DATA  =>  ROM8_DATA22_SIG,
    ROM23_DATA  =>  ROM8_DATA23_SIG,
    ROM24_DATA  =>  ROM8_DATA24_SIG,
    ROM25_DATA  =>  ROM8_DATA25_SIG,
    ROM26_DATA  =>  ROM8_DATA26_SIG,
    ROM27_DATA  =>  ROM8_DATA27_SIG,
    ROM28_DATA  =>  ROM8_DATA28_SIG,
    ROM29_DATA  =>  ROM8_DATA29_SIG,
    ADDR0       =>  ADDR8_0_SIG,
    ADDR1       =>  ADDR8_1_SIG,
    ADDR2       =>  ADDR8_2_SIG,
    ADDR3       =>  ADDR8_3_SIG,
    ADDR4       =>  ADDR8_4_SIG,
    ADDR5       =>  ADDR8_5_SIG,
    ADDR6       =>  ADDR8_6_SIG,
    ADDR7       =>  ADDR8_7_SIG,
    ADDR8       =>  ADDR8_8_SIG,
    ADDR9       =>  ADDR8_9_SIG,
    ADDR10      =>  ADDR8_10_SIG,
    ADDR11      =>  ADDR8_11_SIG,
    ADDR12      =>  ADDR8_12_SIG,
    ADDR13      =>  ADDR8_13_SIG,
    ADDR14      =>  ADDR8_14_SIG,
    ADDR15      =>  ADDR8_15_SIG,
    ADDR16      =>  ADDR8_16_SIG,
    ADDR17      =>  ADDR8_17_SIG,
    ADDR18      =>  ADDR8_18_SIG,
    ADDR19      =>  ADDR8_19_SIG,
    ADDR20      =>  ADDR8_20_SIG,
    ADDR21      =>  ADDR8_21_SIG,
    ADDR22      =>  ADDR8_22_SIG,
    ADDR23      =>  ADDR8_23_SIG,
    ADDR24      =>  ADDR8_24_SIG,
    ADDR25      =>  ADDR8_25_SIG,
    ADDR26      =>  ADDR8_26_SIG,
    ADDR27      =>  ADDR8_27_SIG,
    ADDR28      =>  ADDR8_28_SIG,
    ADDR29      =>  ADDR8_29_SIG,
    DOUT        =>  O_VM8_OUT_SIG
);

O_VM9_INST: OUTPUT_VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER => 5)
Port map (
    CLK         =>  CLK,
    RESET       =>  RESET,
    SET         =>  SET_O_VM,
    DIN0        =>  DIN0_SIG,
    DIN1        =>  DIN1_SIG,
    DIN2        =>  DIN2_SIG,
    DIN3        =>  DIN3_SIG,
    DIN4        =>  DIN4_SIG,
    DIN5        =>  DIN5_SIG,
    DIN6        =>  DIN6_SIG,
    DIN7        =>  DIN7_SIG,
    DIN8        =>  DIN8_SIG,
    DIN9        =>  DIN9_SIG,
    DIN10       =>  DIN10_SIG,
    DIN11       =>  DIN11_SIG,
    DIN12       =>  DIN12_SIG,
    DIN13       =>  DIN13_SIG,
    DIN14       =>  DIN14_SIG,
    DIN15       =>  DIN15_SIG,
    DIN16       =>  DIN16_SIG,
    DIN17       =>  DIN17_SIG,
    DIN18       =>  DIN18_SIG,
    DIN19       =>  DIN19_SIG,
    DIN20       =>  DIN20_SIG,
    DIN21       =>  DIN21_SIG,
    DIN22       =>  DIN22_SIG,
    DIN23       =>  DIN23_SIG,
    DIN24       =>  DIN24_SIG,
    DIN25       =>  DIN25_SIG,
    DIN26       =>  DIN26_SIG,
    DIN27       =>  DIN27_SIG,
    DIN28       =>  DIN28_SIG,
    DIN29       =>  DIN29_SIG,
    ROM0_DATA   =>  ROM9_DATA0_SIG,
    ROM1_DATA   =>  ROM9_DATA1_SIG,
    ROM2_DATA   =>  ROM9_DATA2_SIG,
    ROM3_DATA   =>  ROM9_DATA3_SIG,
    ROM4_DATA   =>  ROM9_DATA4_SIG,
    ROM5_DATA   =>  ROM9_DATA5_SIG,
    ROM6_DATA   =>  ROM9_DATA6_SIG,
    ROM7_DATA   =>  ROM9_DATA7_SIG,
    ROM8_DATA   =>  ROM9_DATA8_SIG,
    ROM9_DATA   =>  ROM9_DATA9_SIG,
    ROM10_DATA  =>  ROM9_DATA10_SIG,
    ROM11_DATA  =>  ROM9_DATA11_SIG,
    ROM12_DATA  =>  ROM9_DATA12_SIG,
    ROM13_DATA  =>  ROM9_DATA13_SIG,
    ROM14_DATA  =>  ROM9_DATA14_SIG,
    ROM15_DATA  =>  ROM9_DATA15_SIG,
    ROM16_DATA  =>  ROM9_DATA16_SIG,
    ROM17_DATA  =>  ROM9_DATA17_SIG,
    ROM18_DATA  =>  ROM9_DATA18_SIG,
    ROM19_DATA  =>  ROM9_DATA19_SIG,
    ROM20_DATA  =>  ROM9_DATA20_SIG,
    ROM21_DATA  =>  ROM9_DATA21_SIG,
    ROM22_DATA  =>  ROM9_DATA22_SIG,
    ROM23_DATA  =>  ROM9_DATA23_SIG,
    ROM24_DATA  =>  ROM9_DATA24_SIG,
    ROM25_DATA  =>  ROM9_DATA25_SIG,
    ROM26_DATA  =>  ROM9_DATA26_SIG,
    ROM27_DATA  =>  ROM9_DATA27_SIG,
    ROM28_DATA  =>  ROM9_DATA28_SIG,
    ROM29_DATA  =>  ROM9_DATA29_SIG,
    ADDR0       =>  ADDR9_0_SIG,
    ADDR1       =>  ADDR9_1_SIG,
    ADDR2       =>  ADDR9_2_SIG,
    ADDR3       =>  ADDR9_3_SIG,
    ADDR4       =>  ADDR9_4_SIG,
    ADDR5       =>  ADDR9_5_SIG,
    ADDR6       =>  ADDR9_6_SIG,
    ADDR7       =>  ADDR9_7_SIG,
    ADDR8       =>  ADDR9_8_SIG,
    ADDR9       =>  ADDR9_9_SIG,
    ADDR10      =>  ADDR9_10_SIG,
    ADDR11      =>  ADDR9_11_SIG,
    ADDR12      =>  ADDR9_12_SIG,
    ADDR13      =>  ADDR9_13_SIG,
    ADDR14      =>  ADDR9_14_SIG,
    ADDR15      =>  ADDR9_15_SIG,
    ADDR16      =>  ADDR9_16_SIG,
    ADDR17      =>  ADDR9_17_SIG,
    ADDR18      =>  ADDR9_18_SIG,
    ADDR19      =>  ADDR9_19_SIG,
    ADDR20      =>  ADDR9_20_SIG,
    ADDR21      =>  ADDR9_21_SIG,
    ADDR22      =>  ADDR9_22_SIG,
    ADDR23      =>  ADDR9_23_SIG,
    ADDR24      =>  ADDR9_24_SIG,
    ADDR25      =>  ADDR9_25_SIG,
    ADDR26      =>  ADDR9_26_SIG,
    ADDR27      =>  ADDR9_27_SIG,
    ADDR28      =>  ADDR9_28_SIG,
    ADDR29      =>  ADDR9_29_SIG,
    DOUT        =>  O_VM9_OUT_SIG
);

OUTPUT_WEIGHT_ROM0_INST: OUTPUT_WEIGHT_ROM
Generic map( WIDTH => 32,
             POWER => 5 ) 
Port map ( 
    ADDR0  => ADDR0_0_SIG,
    ADDR1  => ADDR0_1_SIG,
    ADDR2  => ADDR0_2_SIG,
    ADDR3  => ADDR0_3_SIG,
    ADDR4  => ADDR0_4_SIG,
    ADDR5  => ADDR0_5_SIG,
    ADDR6  => ADDR0_6_SIG,
    ADDR7  => ADDR0_7_SIG,
    ADDR8  => ADDR0_8_SIG,
    ADDR9  => ADDR0_9_SIG,
    ADDR10 => ADDR0_10_SIG,
    ADDR11 => ADDR0_11_SIG,
    ADDR12 => ADDR0_12_SIG,
    ADDR13 => ADDR0_13_SIG,
    ADDR14 => ADDR0_14_SIG,
    ADDR15 => ADDR0_15_SIG,
    ADDR16 => ADDR0_16_SIG,
    ADDR17 => ADDR0_17_SIG,
    ADDR18 => ADDR0_18_SIG,
    ADDR19 => ADDR0_19_SIG,
    ADDR20 => ADDR0_20_SIG,
    ADDR21 => ADDR0_21_SIG,
    ADDR22 => ADDR0_22_SIG,
    ADDR23 => ADDR0_23_SIG,
    ADDR24 => ADDR0_24_SIG,
    ADDR25 => ADDR0_25_SIG,
    ADDR26 => ADDR0_26_SIG,
    ADDR27 => ADDR0_27_SIG,
    ADDR28 => ADDR0_28_SIG,
    ADDR29 => ADDR0_29_SIG,
    DATA0  => ROM0_DATA0_SIG,
    DATA1  => ROM0_DATA1_SIG,
    DATA2  => ROM0_DATA2_SIG,
    DATA3  => ROM0_DATA3_SIG,
    DATA4  => ROM0_DATA4_SIG,
    DATA5  => ROM0_DATA5_SIG,
    DATA6  => ROM0_DATA6_SIG,
    DATA7  => ROM0_DATA7_SIG,
    DATA8  => ROM0_DATA8_SIG,
    DATA9  => ROM0_DATA9_SIG,
    DATA10 => ROM0_DATA10_SIG,
    DATA11 => ROM0_DATA11_SIG,
    DATA12 => ROM0_DATA12_SIG,
    DATA13 => ROM0_DATA13_SIG,
    DATA14 => ROM0_DATA14_SIG,
    DATA15 => ROM0_DATA15_SIG,
    DATA16 => ROM0_DATA16_SIG,
    DATA17 => ROM0_DATA17_SIG,
    DATA18 => ROM0_DATA18_SIG,
    DATA19 => ROM0_DATA19_SIG,
    DATA20 => ROM0_DATA20_SIG,
    DATA21 => ROM0_DATA21_SIG,
    DATA22 => ROM0_DATA22_SIG,
    DATA23 => ROM0_DATA23_SIG,
    DATA24 => ROM0_DATA24_SIG,
    DATA25 => ROM0_DATA25_SIG,
    DATA26 => ROM0_DATA26_SIG,
    DATA27 => ROM0_DATA27_SIG,
    DATA28 => ROM0_DATA28_SIG,
    DATA29 => ROM0_DATA29_SIG
);

OUTPUT_WEIGHT_ROM1_INST: OUTPUT_WEIGHT_ROM
Generic map( WIDTH => 32,
             POWER => 5 ) 
Port map ( 
    ADDR0  => ADDR1_0_SIG,
    ADDR1  => ADDR1_1_SIG,
    ADDR2  => ADDR1_2_SIG,
    ADDR3  => ADDR1_3_SIG,
    ADDR4  => ADDR1_4_SIG,
    ADDR5  => ADDR1_5_SIG,
    ADDR6  => ADDR1_6_SIG,
    ADDR7  => ADDR1_7_SIG,
    ADDR8  => ADDR1_8_SIG,
    ADDR9  => ADDR1_9_SIG,
    ADDR10 => ADDR1_10_SIG,
    ADDR11 => ADDR1_11_SIG,
    ADDR12 => ADDR1_12_SIG,
    ADDR13 => ADDR1_13_SIG,
    ADDR14 => ADDR1_14_SIG,
    ADDR15 => ADDR1_15_SIG,
    ADDR16 => ADDR1_16_SIG,
    ADDR17 => ADDR1_17_SIG,
    ADDR18 => ADDR1_18_SIG,
    ADDR19 => ADDR1_19_SIG,
    ADDR20 => ADDR1_20_SIG,
    ADDR21 => ADDR1_21_SIG,
    ADDR22 => ADDR1_22_SIG,
    ADDR23 => ADDR1_23_SIG,
    ADDR24 => ADDR1_24_SIG,
    ADDR25 => ADDR1_25_SIG,
    ADDR26 => ADDR1_26_SIG,
    ADDR27 => ADDR1_27_SIG,
    ADDR28 => ADDR1_28_SIG,
    ADDR29 => ADDR1_29_SIG,
    DATA0  => ROM1_DATA0_SIG,
    DATA1  => ROM1_DATA1_SIG,
    DATA2  => ROM1_DATA2_SIG,
    DATA3  => ROM1_DATA3_SIG,
    DATA4  => ROM1_DATA4_SIG,
    DATA5  => ROM1_DATA5_SIG,
    DATA6  => ROM1_DATA6_SIG,
    DATA7  => ROM1_DATA7_SIG,
    DATA8  => ROM1_DATA8_SIG,
    DATA9  => ROM1_DATA9_SIG,
    DATA10 => ROM1_DATA10_SIG,
    DATA11 => ROM1_DATA11_SIG,
    DATA12 => ROM1_DATA12_SIG,
    DATA13 => ROM1_DATA13_SIG,
    DATA14 => ROM1_DATA14_SIG,
    DATA15 => ROM1_DATA15_SIG,
    DATA16 => ROM1_DATA16_SIG,
    DATA17 => ROM1_DATA17_SIG,
    DATA18 => ROM1_DATA18_SIG,
    DATA19 => ROM1_DATA19_SIG,
    DATA20 => ROM1_DATA20_SIG,
    DATA21 => ROM1_DATA21_SIG,
    DATA22 => ROM1_DATA22_SIG,
    DATA23 => ROM1_DATA23_SIG,
    DATA24 => ROM1_DATA24_SIG,
    DATA25 => ROM1_DATA25_SIG,
    DATA26 => ROM1_DATA26_SIG,
    DATA27 => ROM1_DATA27_SIG,
    DATA28 => ROM1_DATA28_SIG,
    DATA29 => ROM1_DATA29_SIG
);

OUTPUT_WEIGHT_ROM2_INST: OUTPUT_WEIGHT_ROM
Generic map( WIDTH => 32,
             POWER => 5 ) 
Port map ( 
    ADDR0  => ADDR2_0_SIG,
    ADDR1  => ADDR2_1_SIG,
    ADDR2  => ADDR2_2_SIG,
    ADDR3  => ADDR2_3_SIG,
    ADDR4  => ADDR2_4_SIG,
    ADDR5  => ADDR2_5_SIG,
    ADDR6  => ADDR2_6_SIG,
    ADDR7  => ADDR2_7_SIG,
    ADDR8  => ADDR2_8_SIG,
    ADDR9  => ADDR2_9_SIG,
    ADDR10 => ADDR2_10_SIG,
    ADDR11 => ADDR2_11_SIG,
    ADDR12 => ADDR2_12_SIG,
    ADDR13 => ADDR2_13_SIG,
    ADDR14 => ADDR2_14_SIG,
    ADDR15 => ADDR2_15_SIG,
    ADDR16 => ADDR2_16_SIG,
    ADDR17 => ADDR2_17_SIG,
    ADDR18 => ADDR2_18_SIG,
    ADDR19 => ADDR2_19_SIG,
    ADDR20 => ADDR2_20_SIG,
    ADDR21 => ADDR2_21_SIG,
    ADDR22 => ADDR2_22_SIG,
    ADDR23 => ADDR2_23_SIG,
    ADDR24 => ADDR2_24_SIG,
    ADDR25 => ADDR2_25_SIG,
    ADDR26 => ADDR2_26_SIG,
    ADDR27 => ADDR2_27_SIG,
    ADDR28 => ADDR2_28_SIG,
    ADDR29 => ADDR2_29_SIG,
    DATA0  => ROM2_DATA0_SIG,
    DATA1  => ROM2_DATA1_SIG,
    DATA2  => ROM2_DATA2_SIG,
    DATA3  => ROM2_DATA3_SIG,
    DATA4  => ROM2_DATA4_SIG,
    DATA5  => ROM2_DATA5_SIG,
    DATA6  => ROM2_DATA6_SIG,
    DATA7  => ROM2_DATA7_SIG,
    DATA8  => ROM2_DATA8_SIG,
    DATA9  => ROM2_DATA9_SIG,
    DATA10 => ROM2_DATA10_SIG,
    DATA11 => ROM2_DATA11_SIG,
    DATA12 => ROM2_DATA12_SIG,
    DATA13 => ROM2_DATA13_SIG,
    DATA14 => ROM2_DATA14_SIG,
    DATA15 => ROM2_DATA15_SIG,
    DATA16 => ROM2_DATA16_SIG,
    DATA17 => ROM2_DATA17_SIG,
    DATA18 => ROM2_DATA18_SIG,
    DATA19 => ROM2_DATA19_SIG,
    DATA20 => ROM2_DATA20_SIG,
    DATA21 => ROM2_DATA21_SIG,
    DATA22 => ROM2_DATA22_SIG,
    DATA23 => ROM2_DATA23_SIG,
    DATA24 => ROM2_DATA24_SIG,
    DATA25 => ROM2_DATA25_SIG,
    DATA26 => ROM2_DATA26_SIG,
    DATA27 => ROM2_DATA27_SIG,
    DATA28 => ROM2_DATA28_SIG,
    DATA29 => ROM2_DATA29_SIG
);

OUTPUT_WEIGHT_ROM3_INST: OUTPUT_WEIGHT_ROM
Generic map( WIDTH => 32,
             POWER => 5 ) 
Port map ( 
    ADDR0  => ADDR3_0_SIG,
    ADDR1  => ADDR3_1_SIG,
    ADDR2  => ADDR3_2_SIG,
    ADDR3  => ADDR3_3_SIG,
    ADDR4  => ADDR3_4_SIG,
    ADDR5  => ADDR3_5_SIG,
    ADDR6  => ADDR3_6_SIG,
    ADDR7  => ADDR3_7_SIG,
    ADDR8  => ADDR3_8_SIG,
    ADDR9  => ADDR3_9_SIG,
    ADDR10 => ADDR3_10_SIG,
    ADDR11 => ADDR3_11_SIG,
    ADDR12 => ADDR3_12_SIG,
    ADDR13 => ADDR3_13_SIG,
    ADDR14 => ADDR3_14_SIG,
    ADDR15 => ADDR3_15_SIG,
    ADDR16 => ADDR3_16_SIG,
    ADDR17 => ADDR3_17_SIG,
    ADDR18 => ADDR3_18_SIG,
    ADDR19 => ADDR3_19_SIG,
    ADDR20 => ADDR3_20_SIG,
    ADDR21 => ADDR3_21_SIG,
    ADDR22 => ADDR3_22_SIG,
    ADDR23 => ADDR3_23_SIG,
    ADDR24 => ADDR3_24_SIG,
    ADDR25 => ADDR3_25_SIG,
    ADDR26 => ADDR3_26_SIG,
    ADDR27 => ADDR3_27_SIG,
    ADDR28 => ADDR3_28_SIG,
    ADDR29 => ADDR3_29_SIG,
    DATA0  => ROM3_DATA0_SIG,
    DATA1  => ROM3_DATA1_SIG,
    DATA2  => ROM3_DATA2_SIG,
    DATA3  => ROM3_DATA3_SIG,
    DATA4  => ROM3_DATA4_SIG,
    DATA5  => ROM3_DATA5_SIG,
    DATA6  => ROM3_DATA6_SIG,
    DATA7  => ROM3_DATA7_SIG,
    DATA8  => ROM3_DATA8_SIG,
    DATA9  => ROM3_DATA9_SIG,
    DATA10 => ROM3_DATA10_SIG,
    DATA11 => ROM3_DATA11_SIG,
    DATA12 => ROM3_DATA12_SIG,
    DATA13 => ROM3_DATA13_SIG,
    DATA14 => ROM3_DATA14_SIG,
    DATA15 => ROM3_DATA15_SIG,
    DATA16 => ROM3_DATA16_SIG,
    DATA17 => ROM3_DATA17_SIG,
    DATA18 => ROM3_DATA18_SIG,
    DATA19 => ROM3_DATA19_SIG,
    DATA20 => ROM3_DATA20_SIG,
    DATA21 => ROM3_DATA21_SIG,
    DATA22 => ROM3_DATA22_SIG,
    DATA23 => ROM3_DATA23_SIG,
    DATA24 => ROM3_DATA24_SIG,
    DATA25 => ROM3_DATA25_SIG,
    DATA26 => ROM3_DATA26_SIG,
    DATA27 => ROM3_DATA27_SIG,
    DATA28 => ROM3_DATA28_SIG,
    DATA29 => ROM3_DATA29_SIG
);

OUTPUT_WEIGHT_ROM4_INST: OUTPUT_WEIGHT_ROM
Generic map( WIDTH => 32,
             POWER => 5 ) 
Port map ( 
    ADDR0  => ADDR4_0_SIG,
    ADDR1  => ADDR4_1_SIG,
    ADDR2  => ADDR4_2_SIG,
    ADDR3  => ADDR4_3_SIG,
    ADDR4  => ADDR4_4_SIG,
    ADDR5  => ADDR4_5_SIG,
    ADDR6  => ADDR4_6_SIG,
    ADDR7  => ADDR4_7_SIG,
    ADDR8  => ADDR4_8_SIG,
    ADDR9  => ADDR4_9_SIG,
    ADDR10 => ADDR4_10_SIG,
    ADDR11 => ADDR4_11_SIG,
    ADDR12 => ADDR4_12_SIG,
    ADDR13 => ADDR4_13_SIG,
    ADDR14 => ADDR4_14_SIG,
    ADDR15 => ADDR4_15_SIG,
    ADDR16 => ADDR4_16_SIG,
    ADDR17 => ADDR4_17_SIG,
    ADDR18 => ADDR4_18_SIG,
    ADDR19 => ADDR4_19_SIG,
    ADDR20 => ADDR4_20_SIG,
    ADDR21 => ADDR4_21_SIG,
    ADDR22 => ADDR4_22_SIG,
    ADDR23 => ADDR4_23_SIG,
    ADDR24 => ADDR4_24_SIG,
    ADDR25 => ADDR4_25_SIG,
    ADDR26 => ADDR4_26_SIG,
    ADDR27 => ADDR4_27_SIG,
    ADDR28 => ADDR4_28_SIG,
    ADDR29 => ADDR4_29_SIG,
    DATA0  => ROM4_DATA0_SIG,
    DATA1  => ROM4_DATA1_SIG,
    DATA2  => ROM4_DATA2_SIG,
    DATA3  => ROM4_DATA3_SIG,
    DATA4  => ROM4_DATA4_SIG,
    DATA5  => ROM4_DATA5_SIG,
    DATA6  => ROM4_DATA6_SIG,
    DATA7  => ROM4_DATA7_SIG,
    DATA8  => ROM4_DATA8_SIG,
    DATA9  => ROM4_DATA9_SIG,
    DATA10 => ROM4_DATA10_SIG,
    DATA11 => ROM4_DATA11_SIG,
    DATA12 => ROM4_DATA12_SIG,
    DATA13 => ROM4_DATA13_SIG,
    DATA14 => ROM4_DATA14_SIG,
    DATA15 => ROM4_DATA15_SIG,
    DATA16 => ROM4_DATA16_SIG,
    DATA17 => ROM4_DATA17_SIG,
    DATA18 => ROM4_DATA18_SIG,
    DATA19 => ROM4_DATA19_SIG,
    DATA20 => ROM4_DATA20_SIG,
    DATA21 => ROM4_DATA21_SIG,
    DATA22 => ROM4_DATA22_SIG,
    DATA23 => ROM4_DATA23_SIG,
    DATA24 => ROM4_DATA24_SIG,
    DATA25 => ROM4_DATA25_SIG,
    DATA26 => ROM4_DATA26_SIG,
    DATA27 => ROM4_DATA27_SIG,
    DATA28 => ROM4_DATA28_SIG,
    DATA29 => ROM4_DATA29_SIG
);

OUTPUT_WEIGHT_ROM5_INST: OUTPUT_WEIGHT_ROM
Generic map( WIDTH => 32,
             POWER => 5 ) 
Port map ( 
    ADDR0  => ADDR5_0_SIG,
    ADDR1  => ADDR5_1_SIG,
    ADDR2  => ADDR5_2_SIG,
    ADDR3  => ADDR5_3_SIG,
    ADDR4  => ADDR5_4_SIG,
    ADDR5  => ADDR5_5_SIG,
    ADDR6  => ADDR5_6_SIG,
    ADDR7  => ADDR5_7_SIG,
    ADDR8  => ADDR5_8_SIG,
    ADDR9  => ADDR5_9_SIG,
    ADDR10 => ADDR5_10_SIG,
    ADDR11 => ADDR5_11_SIG,
    ADDR12 => ADDR5_12_SIG,
    ADDR13 => ADDR5_13_SIG,
    ADDR14 => ADDR5_14_SIG,
    ADDR15 => ADDR5_15_SIG,
    ADDR16 => ADDR5_16_SIG,
    ADDR17 => ADDR5_17_SIG,
    ADDR18 => ADDR5_18_SIG,
    ADDR19 => ADDR5_19_SIG,
    ADDR20 => ADDR5_20_SIG,
    ADDR21 => ADDR5_21_SIG,
    ADDR22 => ADDR5_22_SIG,
    ADDR23 => ADDR5_23_SIG,
    ADDR24 => ADDR5_24_SIG,
    ADDR25 => ADDR5_25_SIG,
    ADDR26 => ADDR5_26_SIG,
    ADDR27 => ADDR5_27_SIG,
    ADDR28 => ADDR5_28_SIG,
    ADDR29 => ADDR5_29_SIG,
    DATA0  => ROM5_DATA0_SIG,
    DATA1  => ROM5_DATA1_SIG,
    DATA2  => ROM5_DATA2_SIG,
    DATA3  => ROM5_DATA3_SIG,
    DATA4  => ROM5_DATA4_SIG,
    DATA5  => ROM5_DATA5_SIG,
    DATA6  => ROM5_DATA6_SIG,
    DATA7  => ROM5_DATA7_SIG,
    DATA8  => ROM5_DATA8_SIG,
    DATA9  => ROM5_DATA9_SIG,
    DATA10 => ROM5_DATA10_SIG,
    DATA11 => ROM5_DATA11_SIG,
    DATA12 => ROM5_DATA12_SIG,
    DATA13 => ROM5_DATA13_SIG,
    DATA14 => ROM5_DATA14_SIG,
    DATA15 => ROM5_DATA15_SIG,
    DATA16 => ROM5_DATA16_SIG,
    DATA17 => ROM5_DATA17_SIG,
    DATA18 => ROM5_DATA18_SIG,
    DATA19 => ROM5_DATA19_SIG,
    DATA20 => ROM5_DATA20_SIG,
    DATA21 => ROM5_DATA21_SIG,
    DATA22 => ROM5_DATA22_SIG,
    DATA23 => ROM5_DATA23_SIG,
    DATA24 => ROM5_DATA24_SIG,
    DATA25 => ROM5_DATA25_SIG,
    DATA26 => ROM5_DATA26_SIG,
    DATA27 => ROM5_DATA27_SIG,
    DATA28 => ROM5_DATA28_SIG,
    DATA29 => ROM5_DATA29_SIG
);

OUTPUT_WEIGHT_ROM6_INST: OUTPUT_WEIGHT_ROM
Generic map( WIDTH => 32,
             POWER => 5 ) 
Port map ( 
    ADDR0  => ADDR6_0_SIG,
    ADDR1  => ADDR6_1_SIG,
    ADDR2  => ADDR6_2_SIG,
    ADDR3  => ADDR6_3_SIG,
    ADDR4  => ADDR6_4_SIG,
    ADDR5  => ADDR6_5_SIG,
    ADDR6  => ADDR6_6_SIG,
    ADDR7  => ADDR6_7_SIG,
    ADDR8  => ADDR6_8_SIG,
    ADDR9  => ADDR6_9_SIG,
    ADDR10 => ADDR6_10_SIG,
    ADDR11 => ADDR6_11_SIG,
    ADDR12 => ADDR6_12_SIG,
    ADDR13 => ADDR6_13_SIG,
    ADDR14 => ADDR6_14_SIG,
    ADDR15 => ADDR6_15_SIG,
    ADDR16 => ADDR6_16_SIG,
    ADDR17 => ADDR6_17_SIG,
    ADDR18 => ADDR6_18_SIG,
    ADDR19 => ADDR6_19_SIG,
    ADDR20 => ADDR6_20_SIG,
    ADDR21 => ADDR6_21_SIG,
    ADDR22 => ADDR6_22_SIG,
    ADDR23 => ADDR6_23_SIG,
    ADDR24 => ADDR6_24_SIG,
    ADDR25 => ADDR6_25_SIG,
    ADDR26 => ADDR6_26_SIG,
    ADDR27 => ADDR6_27_SIG,
    ADDR28 => ADDR6_28_SIG,
    ADDR29 => ADDR6_29_SIG,
    DATA0  => ROM6_DATA0_SIG,
    DATA1  => ROM6_DATA1_SIG,
    DATA2  => ROM6_DATA2_SIG,
    DATA3  => ROM6_DATA3_SIG,
    DATA4  => ROM6_DATA4_SIG,
    DATA5  => ROM6_DATA5_SIG,
    DATA6  => ROM6_DATA6_SIG,
    DATA7  => ROM6_DATA7_SIG,
    DATA8  => ROM6_DATA8_SIG,
    DATA9  => ROM6_DATA9_SIG,
    DATA10 => ROM6_DATA10_SIG,
    DATA11 => ROM6_DATA11_SIG,
    DATA12 => ROM6_DATA12_SIG,
    DATA13 => ROM6_DATA13_SIG,
    DATA14 => ROM6_DATA14_SIG,
    DATA15 => ROM6_DATA15_SIG,
    DATA16 => ROM6_DATA16_SIG,
    DATA17 => ROM6_DATA17_SIG,
    DATA18 => ROM6_DATA18_SIG,
    DATA19 => ROM6_DATA19_SIG,
    DATA20 => ROM6_DATA20_SIG,
    DATA21 => ROM6_DATA21_SIG,
    DATA22 => ROM6_DATA22_SIG,
    DATA23 => ROM6_DATA23_SIG,
    DATA24 => ROM6_DATA24_SIG,
    DATA25 => ROM6_DATA25_SIG,
    DATA26 => ROM6_DATA26_SIG,
    DATA27 => ROM6_DATA27_SIG,
    DATA28 => ROM6_DATA28_SIG,
    DATA29 => ROM6_DATA29_SIG
);

OUTPUT_WEIGHT_ROM7_INST: OUTPUT_WEIGHT_ROM
Generic map( WIDTH => 32,
             POWER => 5 ) 
Port map ( 
    ADDR0  => ADDR7_0_SIG,
    ADDR1  => ADDR7_1_SIG,
    ADDR2  => ADDR7_2_SIG,
    ADDR3  => ADDR7_3_SIG,
    ADDR4  => ADDR7_4_SIG,
    ADDR5  => ADDR7_5_SIG,
    ADDR6  => ADDR7_6_SIG,
    ADDR7  => ADDR7_7_SIG,
    ADDR8  => ADDR7_8_SIG,
    ADDR9  => ADDR7_9_SIG,
    ADDR10 => ADDR7_10_SIG,
    ADDR11 => ADDR7_11_SIG,
    ADDR12 => ADDR7_12_SIG,
    ADDR13 => ADDR7_13_SIG,
    ADDR14 => ADDR7_14_SIG,
    ADDR15 => ADDR7_15_SIG,
    ADDR16 => ADDR7_16_SIG,
    ADDR17 => ADDR7_17_SIG,
    ADDR18 => ADDR7_18_SIG,
    ADDR19 => ADDR7_19_SIG,
    ADDR20 => ADDR7_20_SIG,
    ADDR21 => ADDR7_21_SIG,
    ADDR22 => ADDR7_22_SIG,
    ADDR23 => ADDR7_23_SIG,
    ADDR24 => ADDR7_24_SIG,
    ADDR25 => ADDR7_25_SIG,
    ADDR26 => ADDR7_26_SIG,
    ADDR27 => ADDR7_27_SIG,
    ADDR28 => ADDR7_28_SIG,
    ADDR29 => ADDR7_29_SIG,
    DATA0  => ROM7_DATA0_SIG,
    DATA1  => ROM7_DATA1_SIG,
    DATA2  => ROM7_DATA2_SIG,
    DATA3  => ROM7_DATA3_SIG,
    DATA4  => ROM7_DATA4_SIG,
    DATA5  => ROM7_DATA5_SIG,
    DATA6  => ROM7_DATA6_SIG,
    DATA7  => ROM7_DATA7_SIG,
    DATA8  => ROM7_DATA8_SIG,
    DATA9  => ROM7_DATA9_SIG,
    DATA10 => ROM7_DATA10_SIG,
    DATA11 => ROM7_DATA11_SIG,
    DATA12 => ROM7_DATA12_SIG,
    DATA13 => ROM7_DATA13_SIG,
    DATA14 => ROM7_DATA14_SIG,
    DATA15 => ROM7_DATA15_SIG,
    DATA16 => ROM7_DATA16_SIG,
    DATA17 => ROM7_DATA17_SIG,
    DATA18 => ROM7_DATA18_SIG,
    DATA19 => ROM7_DATA19_SIG,
    DATA20 => ROM7_DATA20_SIG,
    DATA21 => ROM7_DATA21_SIG,
    DATA22 => ROM7_DATA22_SIG,
    DATA23 => ROM7_DATA23_SIG,
    DATA24 => ROM7_DATA24_SIG,
    DATA25 => ROM7_DATA25_SIG,
    DATA26 => ROM7_DATA26_SIG,
    DATA27 => ROM7_DATA27_SIG,
    DATA28 => ROM7_DATA28_SIG,
    DATA29 => ROM7_DATA29_SIG
);

OUTPUT_WEIGHT_ROM8_INST: OUTPUT_WEIGHT_ROM
Generic map( WIDTH => 32,
             POWER => 5 ) 
Port map ( 
    ADDR0  => ADDR8_0_SIG,
    ADDR1  => ADDR8_1_SIG,
    ADDR2  => ADDR8_2_SIG,
    ADDR3  => ADDR8_3_SIG,
    ADDR4  => ADDR8_4_SIG,
    ADDR5  => ADDR8_5_SIG,
    ADDR6  => ADDR8_6_SIG,
    ADDR7  => ADDR8_7_SIG,
    ADDR8  => ADDR8_8_SIG,
    ADDR9  => ADDR8_9_SIG,
    ADDR10 => ADDR8_10_SIG,
    ADDR11 => ADDR8_11_SIG,
    ADDR12 => ADDR8_12_SIG,
    ADDR13 => ADDR8_13_SIG,
    ADDR14 => ADDR8_14_SIG,
    ADDR15 => ADDR8_15_SIG,
    ADDR16 => ADDR8_16_SIG,
    ADDR17 => ADDR8_17_SIG,
    ADDR18 => ADDR8_18_SIG,
    ADDR19 => ADDR8_19_SIG,
    ADDR20 => ADDR8_20_SIG,
    ADDR21 => ADDR8_21_SIG,
    ADDR22 => ADDR8_22_SIG,
    ADDR23 => ADDR8_23_SIG,
    ADDR24 => ADDR8_24_SIG,
    ADDR25 => ADDR8_25_SIG,
    ADDR26 => ADDR8_26_SIG,
    ADDR27 => ADDR8_27_SIG,
    ADDR28 => ADDR8_28_SIG,
    ADDR29 => ADDR8_29_SIG,
    DATA0  => ROM8_DATA0_SIG,
    DATA1  => ROM8_DATA1_SIG,
    DATA2  => ROM8_DATA2_SIG,
    DATA3  => ROM8_DATA3_SIG,
    DATA4  => ROM8_DATA4_SIG,
    DATA5  => ROM8_DATA5_SIG,
    DATA6  => ROM8_DATA6_SIG,
    DATA7  => ROM8_DATA7_SIG,
    DATA8  => ROM8_DATA8_SIG,
    DATA9  => ROM8_DATA9_SIG,
    DATA10 => ROM8_DATA10_SIG,
    DATA11 => ROM8_DATA11_SIG,
    DATA12 => ROM8_DATA12_SIG,
    DATA13 => ROM8_DATA13_SIG,
    DATA14 => ROM8_DATA14_SIG,
    DATA15 => ROM8_DATA15_SIG,
    DATA16 => ROM8_DATA16_SIG,
    DATA17 => ROM8_DATA17_SIG,
    DATA18 => ROM8_DATA18_SIG,
    DATA19 => ROM8_DATA19_SIG,
    DATA20 => ROM8_DATA20_SIG,
    DATA21 => ROM8_DATA21_SIG,
    DATA22 => ROM8_DATA22_SIG,
    DATA23 => ROM8_DATA23_SIG,
    DATA24 => ROM8_DATA24_SIG,
    DATA25 => ROM8_DATA25_SIG,
    DATA26 => ROM8_DATA26_SIG,
    DATA27 => ROM8_DATA27_SIG,
    DATA28 => ROM8_DATA28_SIG,
    DATA29 => ROM8_DATA29_SIG
);

OUTPUT_WEIGHT_ROM9_INST: OUTPUT_WEIGHT_ROM
Generic map( WIDTH => 32,
             POWER => 5 ) 
Port map ( 
    ADDR0  => ADDR9_0_SIG,
    ADDR1  => ADDR9_1_SIG,
    ADDR2  => ADDR9_2_SIG,
    ADDR3  => ADDR9_3_SIG,
    ADDR4  => ADDR9_4_SIG,
    ADDR5  => ADDR9_5_SIG,
    ADDR6  => ADDR9_6_SIG,
    ADDR7  => ADDR9_7_SIG,
    ADDR8  => ADDR9_8_SIG,
    ADDR9  => ADDR9_9_SIG,
    ADDR10 => ADDR9_10_SIG,
    ADDR11 => ADDR9_11_SIG,
    ADDR12 => ADDR9_12_SIG,
    ADDR13 => ADDR9_13_SIG,
    ADDR14 => ADDR9_14_SIG,
    ADDR15 => ADDR9_15_SIG,
    ADDR16 => ADDR9_16_SIG,
    ADDR17 => ADDR9_17_SIG,
    ADDR18 => ADDR9_18_SIG,
    ADDR19 => ADDR9_19_SIG,
    ADDR20 => ADDR9_20_SIG,
    ADDR21 => ADDR9_21_SIG,
    ADDR22 => ADDR9_22_SIG,
    ADDR23 => ADDR9_23_SIG,
    ADDR24 => ADDR9_24_SIG,
    ADDR25 => ADDR9_25_SIG,
    ADDR26 => ADDR9_26_SIG,
    ADDR27 => ADDR9_27_SIG,
    ADDR28 => ADDR9_28_SIG,
    ADDR29 => ADDR9_29_SIG,
    DATA0  => ROM9_DATA0_SIG,
    DATA1  => ROM9_DATA1_SIG,
    DATA2  => ROM9_DATA2_SIG,
    DATA3  => ROM9_DATA3_SIG,
    DATA4  => ROM9_DATA4_SIG,
    DATA5  => ROM9_DATA5_SIG,
    DATA6  => ROM9_DATA6_SIG,
    DATA7  => ROM9_DATA7_SIG,
    DATA8  => ROM9_DATA8_SIG,
    DATA9  => ROM9_DATA9_SIG,
    DATA10 => ROM9_DATA10_SIG,
    DATA11 => ROM9_DATA11_SIG,
    DATA12 => ROM9_DATA12_SIG,
    DATA13 => ROM9_DATA13_SIG,
    DATA14 => ROM9_DATA14_SIG,
    DATA15 => ROM9_DATA15_SIG,
    DATA16 => ROM9_DATA16_SIG,
    DATA17 => ROM9_DATA17_SIG,
    DATA18 => ROM9_DATA18_SIG,
    DATA19 => ROM9_DATA19_SIG,
    DATA20 => ROM9_DATA20_SIG,
    DATA21 => ROM9_DATA21_SIG,
    DATA22 => ROM9_DATA22_SIG,
    DATA23 => ROM9_DATA23_SIG,
    DATA24 => ROM9_DATA24_SIG,
    DATA25 => ROM9_DATA25_SIG,
    DATA26 => ROM9_DATA26_SIG,
    DATA27 => ROM9_DATA27_SIG,
    DATA28 => ROM9_DATA28_SIG,
    DATA29 => ROM9_DATA29_SIG
);

OUTPUT_BIAS_ROM_INST: OUTPUT_BIAS_ROM
Generic map ( WIDTH => 64,
              POWER => 4) 
Port map ( 
    ADDR0  => BIAS_ADDR0_SIG,
    ADDR1  => BIAS_ADDR1_SIG,
    ADDR2  => BIAS_ADDR2_SIG,
    ADDR3  => BIAS_ADDR3_SIG,
    ADDR4  => BIAS_ADDR4_SIG,
    ADDR5  => BIAS_ADDR5_SIG,
    ADDR6  => BIAS_ADDR6_SIG,
    ADDR7  => BIAS_ADDR7_SIG,
    ADDR8  => BIAS_ADDR8_SIG,
    ADDR9  => BIAS_ADDR9_SIG,
    DATA0  => BIAS0_SIG,
    DATA1  => BIAS1_SIG,
    DATA2  => BIAS2_SIG,
    DATA3  => BIAS3_SIG,
    DATA4  => BIAS4_SIG,
    DATA5  => BIAS5_SIG,
    DATA6  => BIAS6_SIG,
    DATA7  => BIAS7_SIG,
    DATA8  => BIAS8_SIG,
    DATA9  => BIAS9_SIG
);

ADDER0_INST: ADDER
Generic map ( WIDTH => 64)
Port map(
    A    => BIAS0_SIG,
    B    => O_VM0_OUT_SIG,
    S    => ADDER0_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER1_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS1_SIG,
    B    => O_VM1_OUT_SIG,
    S    => ADDER1_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER2_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS2_SIG,
    B    => O_VM2_OUT_SIG,
    S    => ADDER2_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER3_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS3_SIG,
    B    => O_VM3_OUT_SIG,
    S    => ADDER3_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER4_INST: ADDER
Generic map ( WIDTH => 64)
Port map(
    A    => BIAS4_SIG,
    B    => O_VM4_OUT_SIG,
    S    => ADDER4_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER5_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS5_SIG,
    B    => O_VM5_OUT_SIG,
    S    => ADDER5_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER6_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS6_SIG,
    B    => O_VM6_OUT_SIG,
    S    => ADDER6_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER7_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS7_SIG,
    B    => O_VM7_OUT_SIG,
    S    => ADDER7_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER8_INST: ADDER
Generic map ( WIDTH => 64)
Port map(
    A    => BIAS8_SIG,
    B    => O_VM8_OUT_SIG,
    S    => ADDER8_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER9_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS9_SIG,
    B    => O_VM9_OUT_SIG,
    S    => ADDER9_OUT_SIG,
    COUT => open,
    OV   => open
);

RELU_MUX0_INST: RELU_MUX
Generic map ( WIDTH => 64)
Port map (
    DIN  => ADDER0_OUT_SIG,
    DOUT => DOUT0
);

RELU_MUX1_INST: RELU_MUX
Generic map ( WIDTH => 64)
Port map (
    DIN  => ADDER1_OUT_SIG,
    DOUT => DOUT1
);

RELU_MUX2_INST: RELU_MUX
Generic map ( WIDTH => 64)
Port map (
    DIN  => ADDER2_OUT_SIG,
    DOUT => DOUT2
);

RELU_MUX3_INST: RELU_MUX
Generic map ( WIDTH => 64)
Port map (
    DIN  => ADDER3_OUT_SIG,
    DOUT => DOUT3
);

RELU_MUX4_INST: RELU_MUX
Generic map ( WIDTH => 64)
Port map (
    DIN  => ADDER4_OUT_SIG,
    DOUT => DOUT4
);

RELU_MUX5_INST: RELU_MUX
Generic map ( WIDTH => 64)
Port map (
    DIN  => ADDER5_OUT_SIG,
    DOUT => DOUT5
);

RELU_MUX6_INST: RELU_MUX
Generic map ( WIDTH => 64)
Port map (
    DIN  => ADDER6_OUT_SIG,
    DOUT => DOUT6
);

RELU_MUX7_INST: RELU_MUX
Generic map ( WIDTH => 64)
Port map (
    DIN  => ADDER7_OUT_SIG,
    DOUT => DOUT7
);

RELU_MUX8_INST: RELU_MUX
Generic map ( WIDTH => 64)
Port map (
    DIN  => ADDER8_OUT_SIG,
    DOUT => DOUT8
);

RELU_MUX9_INST: RELU_MUX
Generic map ( WIDTH => 64)
Port map (
    DIN  => ADDER9_OUT_SIG,
    DOUT => DOUT9
);

end Structural;
