library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;
--library UNISIM;
--use UNISIM.VComponents.all;

entity FULLY_CONNECTED_LAYER is
Generic (WIDTH : positive := 32;
         POWER : positive := 13);
Port (
    CLK     :  in  std_logic;
    RESET   :  in  std_logic;
    SET_CNT : in  std_logic;
    DIN0    :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN1    :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN2    :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN3    :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN4    :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN5    :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN6    :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN7    :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN8    :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN9    :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN10   :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN11   :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN12   :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN13   :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN14   :   in  std_logic_vector(WIDTH-1 downto 0);
    DIN15   :   in  std_logic_vector(WIDTH-1 downto 0);
    DIN16   :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN17   :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN18   :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN19   :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN20   :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN21   :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN22   :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN23   :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN24   :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN25   :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN26   :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN27   :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN28   :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN29   :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN30   :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN31   :  in  std_logic_vector(WIDTH-1 downto 0);
    DOUT0   :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT1   :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT2   :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT3   :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT4   :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT5   :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT6   :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT7   :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT8   :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT9   :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT10  :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT11  :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT12  :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT13  :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT14  :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT15  :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT16  :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT17  :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT18  :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT19  :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT20  :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT21  :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT22  :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT23  :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT24  :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT25  :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT26  :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT27  :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT28  :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT29  :  out std_logic_vector(WIDTH+WIDTH-1 downto 0);
    SET_CNT_OL : out std_logic
);
end FULLY_CONNECTED_LAYER;

architecture Structural of FULLY_CONNECTED_LAYER is

component VECTOR_MULTIPLIER
Generic(WIDTH : positive := 32;
        POWER : positive := 13);
Port (
    CLK         :  in  std_logic;
    RESET       :  in  std_logic;
    SET         :  in  std_logic;
    DIN0        :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN1        :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN2        :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN3        :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN4        :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN5        :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN6        :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN7        :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN8        :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN9        :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN10       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN11       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN12       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN13       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN14       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN15       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN16       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN17       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN18       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN19       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN20       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN21       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN22       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN23       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN24       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN25       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN26       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN27       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN28       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN29       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN30       :  in  std_logic_vector(WIDTH-1 downto 0);
    DIN31       :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM0_DATA   :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM1_DATA   :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM2_DATA   :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM3_DATA   :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM4_DATA   :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM5_DATA   :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM6_DATA   :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM7_DATA   :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM8_DATA   :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM9_DATA   :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM10_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM11_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM12_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM13_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM14_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM15_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM16_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM17_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM18_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM19_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM20_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM21_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM22_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM23_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM24_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM25_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM26_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM27_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM28_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM29_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM30_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ROM31_DATA  :  in  std_logic_vector(WIDTH-1 downto 0);
    ADDR0       :  out std_logic_vector(POWER-1 downto 0);
    ADDR1       :  out std_logic_vector(POWER-1 downto 0);
    ADDR2       :  out std_logic_vector(POWER-1 downto 0);
    ADDR3       :  out std_logic_vector(POWER-1 downto 0);
    ADDR4       :  out std_logic_vector(POWER-1 downto 0);
    ADDR5       :  out std_logic_vector(POWER-1 downto 0);
    ADDR6       :  out std_logic_vector(POWER-1 downto 0);
    ADDR7       :  out std_logic_vector(POWER-1 downto 0);
    ADDR8       :  out std_logic_vector(POWER-1 downto 0);
    ADDR9       :  out std_logic_vector(POWER-1 downto 0);
    ADDR10      :  out std_logic_vector(POWER-1 downto 0);
    ADDR11      :  out std_logic_vector(POWER-1 downto 0);
    ADDR12      :  out std_logic_vector(POWER-1 downto 0);
    ADDR13      :  out std_logic_vector(POWER-1 downto 0);
    ADDR14      :  out std_logic_vector(POWER-1 downto 0);
    ADDR15      :  out std_logic_vector(POWER-1 downto 0);
    ADDR16      :  out std_logic_vector(POWER-1 downto 0);
    ADDR17      :  out std_logic_vector(POWER-1 downto 0);
    ADDR18      :  out std_logic_vector(POWER-1 downto 0);
    ADDR19      :  out std_logic_vector(POWER-1 downto 0);
    ADDR20      :  out std_logic_vector(POWER-1 downto 0);
    ADDR21      :  out std_logic_vector(POWER-1 downto 0);
    ADDR22      :  out std_logic_vector(POWER-1 downto 0);
    ADDR23      :  out std_logic_vector(POWER-1 downto 0);
    ADDR24      :  out std_logic_vector(POWER-1 downto 0);
    ADDR25      :  out std_logic_vector(POWER-1 downto 0);
    ADDR26      :  out std_logic_vector(POWER-1 downto 0);
    ADDR27      :  out std_logic_vector(POWER-1 downto 0);
    ADDR28      :  out std_logic_vector(POWER-1 downto 0);
    ADDR29      :  out std_logic_vector(POWER-1 downto 0);
    ADDR30      :  out std_logic_vector(POWER-1 downto 0);
    ADDR31      :  out std_logic_vector(POWER-1 downto 0);
    DOUT        :  out std_logic_vector(WIDTH+WIDTH-1 downto 0)
);
end component;

component COUNTER_FOR_FC
Port (
    CLK   :  in  std_logic;
    RESET :  in  std_logic;
    SET   :  in  std_logic;
    COUT1 :  out std_logic;
    COUT2 :  out std_logic
 );
 end component;
 
component WEIGHT_ROM
Generic ( WIDTH : positive := 32;
          POWER : positive := 13); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR26 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR27 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR28 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR29 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR30 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR31 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0);
    DATA26 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA27 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA28 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA29 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA30 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA31 :    out std_logic_vector(WIDTH-1 downto 0)
);
end component; 

component BIAS_ROM_FC
Generic ( WIDTH : positive := 64;
          POWER : positive := 6); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR26 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR27 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR28 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR29 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0);
    DATA26 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA27 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA28 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA29 :    out std_logic_vector(WIDTH-1 downto 0)
);
end component;

component ADDER
Generic ( WIDTH : positive := 32);
Port (
    A    :  in  std_logic_vector(WIDTH-1 downto 0);
    B    :  in  std_logic_vector(WIDTH-1 downto 0);
    S    :  out std_logic_vector(WIDTH-1 downto 0);
    COUT :  out std_logic;
    OV   :  out std_logic
);
end component;

component RELU_MUX
Generic( WIDTH : positive := 32);
Port (
    DIN  :  in  std_logic_vector(WIDTH-1 downto 0);
    DOUT :  out std_logic_vector(WIDTH-1 downto 0)
);
end component;

signal DIN0_SIG, DIN1_SIG, DIN2_SIG, DIN3_SIG, DIN4_SIG, DIN5_SIG, DIN6_SIG, DIN7_SIG,
       DIN8_SIG, DIN9_SIG, DIN10_SIG, DIN11_SIG, DIN12_SIG, DIN13_SIG, DIN14_SIG, DIN15_SIG,
       DIN16_SIG, DIN17_SIG, DIN18_SIG, DIN19_SIG, DIN20_SIG, DIN21_SIG, DIN22_SIG, DIN23_SIG,
       DIN24_SIG, DIN25_SIG, DIN26_SIG, DIN27_SIG, DIN28_SIG, DIN29_SIG, DIN30_SIG, DIN31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM0_DATA0_SIG, ROM0_DATA1_SIG, ROM0_DATA2_SIG, ROM0_DATA3_SIG, ROM0_DATA4_SIG,
       ROM0_DATA5_SIG, ROM0_DATA6_SIG, ROM0_DATA7_SIG, ROM0_DATA8_SIG, ROM0_DATA9_SIG,
       ROM0_DATA10_SIG, ROM0_DATA11_SIG, ROM0_DATA12_SIG, ROM0_DATA13_SIG, ROM0_DATA14_SIG,
       ROM0_DATA15_SIG, ROM0_DATA16_SIG, ROM0_DATA17_SIG, ROM0_DATA18_SIG, ROM0_DATA19_SIG,
       ROM0_DATA20_SIG, ROM0_DATA21_SIG, ROM0_DATA22_SIG, ROM0_DATA23_SIG, ROM0_DATA24_SIG, ROM0_DATA25_SIG,
       ROM0_DATA26_SIG, ROM0_DATA27_SIG, ROM0_DATA28_SIG, ROM0_DATA29_SIG, ROM0_DATA30_SIG, ROM0_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM1_DATA0_SIG, ROM1_DATA1_SIG, ROM1_DATA2_SIG, ROM1_DATA3_SIG, ROM1_DATA4_SIG,
       ROM1_DATA5_SIG, ROM1_DATA6_SIG, ROM1_DATA7_SIG, ROM1_DATA8_SIG, ROM1_DATA9_SIG,
       ROM1_DATA10_SIG, ROM1_DATA11_SIG, ROM1_DATA12_SIG, ROM1_DATA13_SIG, ROM1_DATA14_SIG,
       ROM1_DATA15_SIG, ROM1_DATA16_SIG, ROM1_DATA17_SIG, ROM1_DATA18_SIG, ROM1_DATA19_SIG,
       ROM1_DATA20_SIG, ROM1_DATA21_SIG, ROM1_DATA22_SIG, ROM1_DATA23_SIG, ROM1_DATA24_SIG, ROM1_DATA25_SIG,
       ROM1_DATA26_SIG, ROM1_DATA27_SIG, ROM1_DATA28_SIG, ROM1_DATA29_SIG, ROM1_DATA30_SIG, ROM1_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0'); 
signal ROM2_DATA0_SIG, ROM2_DATA1_SIG, ROM2_DATA2_SIG, ROM2_DATA3_SIG, ROM2_DATA4_SIG,
       ROM2_DATA5_SIG, ROM2_DATA6_SIG, ROM2_DATA7_SIG, ROM2_DATA8_SIG, ROM2_DATA9_SIG,
       ROM2_DATA10_SIG, ROM2_DATA11_SIG, ROM2_DATA12_SIG, ROM2_DATA13_SIG, ROM2_DATA14_SIG,
       ROM2_DATA15_SIG, ROM2_DATA16_SIG, ROM2_DATA17_SIG, ROM2_DATA18_SIG, ROM2_DATA19_SIG,
       ROM2_DATA20_SIG, ROM2_DATA21_SIG, ROM2_DATA22_SIG, ROM2_DATA23_SIG, ROM2_DATA24_SIG, ROM2_DATA25_SIG,
       ROM2_DATA26_SIG, ROM2_DATA27_SIG, ROM2_DATA28_SIG, ROM2_DATA29_SIG, ROM2_DATA30_SIG, ROM2_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM3_DATA0_SIG, ROM3_DATA1_SIG, ROM3_DATA2_SIG, ROM3_DATA3_SIG, ROM3_DATA4_SIG,
       ROM3_DATA5_SIG, ROM3_DATA6_SIG, ROM3_DATA7_SIG, ROM3_DATA8_SIG, ROM3_DATA9_SIG,
       ROM3_DATA10_SIG, ROM3_DATA11_SIG, ROM3_DATA12_SIG, ROM3_DATA13_SIG, ROM3_DATA14_SIG,
       ROM3_DATA15_SIG, ROM3_DATA16_SIG, ROM3_DATA17_SIG, ROM3_DATA18_SIG, ROM3_DATA19_SIG,
       ROM3_DATA20_SIG, ROM3_DATA21_SIG, ROM3_DATA22_SIG, ROM3_DATA23_SIG, ROM3_DATA24_SIG, ROM3_DATA25_SIG,
       ROM3_DATA26_SIG, ROM3_DATA27_SIG, ROM3_DATA28_SIG, ROM3_DATA29_SIG, ROM3_DATA30_SIG, ROM3_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM4_DATA0_SIG, ROM4_DATA1_SIG, ROM4_DATA2_SIG, ROM4_DATA3_SIG, ROM4_DATA4_SIG,
       ROM4_DATA5_SIG, ROM4_DATA6_SIG, ROM4_DATA7_SIG, ROM4_DATA8_SIG, ROM4_DATA9_SIG,
       ROM4_DATA10_SIG, ROM4_DATA11_SIG, ROM4_DATA12_SIG, ROM4_DATA13_SIG, ROM4_DATA14_SIG,
       ROM4_DATA15_SIG, ROM4_DATA16_SIG, ROM4_DATA17_SIG, ROM4_DATA18_SIG, ROM4_DATA19_SIG,
       ROM4_DATA20_SIG, ROM4_DATA21_SIG, ROM4_DATA22_SIG, ROM4_DATA23_SIG, ROM4_DATA24_SIG, ROM4_DATA25_SIG,
       ROM4_DATA26_SIG, ROM4_DATA27_SIG, ROM4_DATA28_SIG, ROM4_DATA29_SIG, ROM4_DATA30_SIG, ROM4_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM5_DATA0_SIG, ROM5_DATA1_SIG, ROM5_DATA2_SIG, ROM5_DATA3_SIG, ROM5_DATA4_SIG,
       ROM5_DATA5_SIG, ROM5_DATA6_SIG, ROM5_DATA7_SIG, ROM5_DATA8_SIG, ROM5_DATA9_SIG,
       ROM5_DATA10_SIG, ROM5_DATA11_SIG, ROM5_DATA12_SIG, ROM5_DATA13_SIG, ROM5_DATA14_SIG,
       ROM5_DATA15_SIG, ROM5_DATA16_SIG, ROM5_DATA17_SIG, ROM5_DATA18_SIG, ROM5_DATA19_SIG,
       ROM5_DATA20_SIG, ROM5_DATA21_SIG, ROM5_DATA22_SIG, ROM5_DATA23_SIG, ROM5_DATA24_SIG, ROM5_DATA25_SIG,
       ROM5_DATA26_SIG, ROM5_DATA27_SIG, ROM5_DATA28_SIG, ROM5_DATA29_SIG, ROM5_DATA30_SIG, ROM5_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM6_DATA0_SIG, ROM6_DATA1_SIG, ROM6_DATA2_SIG, ROM6_DATA3_SIG, ROM6_DATA4_SIG,
       ROM6_DATA5_SIG, ROM6_DATA6_SIG, ROM6_DATA7_SIG, ROM6_DATA8_SIG, ROM6_DATA9_SIG,
       ROM6_DATA10_SIG, ROM6_DATA11_SIG, ROM6_DATA12_SIG, ROM6_DATA13_SIG, ROM6_DATA14_SIG,
       ROM6_DATA15_SIG, ROM6_DATA16_SIG, ROM6_DATA17_SIG, ROM6_DATA18_SIG, ROM6_DATA19_SIG,
       ROM6_DATA20_SIG, ROM6_DATA21_SIG, ROM6_DATA22_SIG, ROM6_DATA23_SIG, ROM6_DATA24_SIG, ROM6_DATA25_SIG,
       ROM6_DATA26_SIG, ROM6_DATA27_SIG, ROM6_DATA28_SIG, ROM6_DATA29_SIG, ROM6_DATA30_SIG, ROM6_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM7_DATA0_SIG, ROM7_DATA1_SIG, ROM7_DATA2_SIG, ROM7_DATA3_SIG, ROM7_DATA4_SIG,
       ROM7_DATA5_SIG, ROM7_DATA6_SIG, ROM7_DATA7_SIG, ROM7_DATA8_SIG, ROM7_DATA9_SIG,
       ROM7_DATA10_SIG, ROM7_DATA11_SIG, ROM7_DATA12_SIG, ROM7_DATA13_SIG, ROM7_DATA14_SIG,
       ROM7_DATA15_SIG, ROM7_DATA16_SIG, ROM7_DATA17_SIG, ROM7_DATA18_SIG, ROM7_DATA19_SIG,
       ROM7_DATA20_SIG, ROM7_DATA21_SIG, ROM7_DATA22_SIG, ROM7_DATA23_SIG, ROM7_DATA24_SIG, ROM7_DATA25_SIG,
       ROM7_DATA26_SIG, ROM7_DATA27_SIG, ROM7_DATA28_SIG, ROM7_DATA29_SIG, ROM7_DATA30_SIG, ROM7_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM8_DATA0_SIG, ROM8_DATA1_SIG, ROM8_DATA2_SIG, ROM8_DATA3_SIG, ROM8_DATA4_SIG,
       ROM8_DATA5_SIG, ROM8_DATA6_SIG, ROM8_DATA7_SIG, ROM8_DATA8_SIG, ROM8_DATA9_SIG,
       ROM8_DATA10_SIG, ROM8_DATA11_SIG, ROM8_DATA12_SIG, ROM8_DATA13_SIG, ROM8_DATA14_SIG,
       ROM8_DATA15_SIG, ROM8_DATA16_SIG, ROM8_DATA17_SIG, ROM8_DATA18_SIG, ROM8_DATA19_SIG,
       ROM8_DATA20_SIG, ROM8_DATA21_SIG, ROM8_DATA22_SIG, ROM8_DATA23_SIG, ROM8_DATA24_SIG, ROM8_DATA25_SIG,
       ROM8_DATA26_SIG, ROM8_DATA27_SIG, ROM8_DATA28_SIG, ROM8_DATA29_SIG, ROM8_DATA30_SIG, ROM8_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM9_DATA0_SIG, ROM9_DATA1_SIG, ROM9_DATA2_SIG, ROM9_DATA3_SIG, ROM9_DATA4_SIG,
       ROM9_DATA5_SIG, ROM9_DATA6_SIG, ROM9_DATA7_SIG, ROM9_DATA8_SIG, ROM9_DATA9_SIG,
       ROM9_DATA10_SIG, ROM9_DATA11_SIG, ROM9_DATA12_SIG, ROM9_DATA13_SIG, ROM9_DATA14_SIG,
       ROM9_DATA15_SIG, ROM9_DATA16_SIG, ROM9_DATA17_SIG, ROM9_DATA18_SIG, ROM9_DATA19_SIG,
       ROM9_DATA20_SIG, ROM9_DATA21_SIG, ROM9_DATA22_SIG, ROM9_DATA23_SIG, ROM9_DATA24_SIG, ROM9_DATA25_SIG,
       ROM9_DATA26_SIG, ROM9_DATA27_SIG, ROM9_DATA28_SIG, ROM9_DATA29_SIG, ROM9_DATA30_SIG, ROM9_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM10_DATA0_SIG, ROM10_DATA1_SIG, ROM10_DATA2_SIG, ROM10_DATA3_SIG, ROM10_DATA4_SIG,
       ROM10_DATA5_SIG, ROM10_DATA6_SIG, ROM10_DATA7_SIG, ROM10_DATA8_SIG, ROM10_DATA9_SIG,
       ROM10_DATA10_SIG, ROM10_DATA11_SIG, ROM10_DATA12_SIG, ROM10_DATA13_SIG, ROM10_DATA14_SIG,
       ROM10_DATA15_SIG, ROM10_DATA16_SIG, ROM10_DATA17_SIG, ROM10_DATA18_SIG, ROM10_DATA19_SIG,
       ROM10_DATA20_SIG, ROM10_DATA21_SIG, ROM10_DATA22_SIG, ROM10_DATA23_SIG, ROM10_DATA24_SIG, ROM10_DATA25_SIG,
       ROM10_DATA26_SIG, ROM10_DATA27_SIG, ROM10_DATA28_SIG, ROM10_DATA29_SIG, ROM10_DATA30_SIG, ROM10_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM11_DATA0_SIG, ROM11_DATA1_SIG, ROM11_DATA2_SIG, ROM11_DATA3_SIG, ROM11_DATA4_SIG,
       ROM11_DATA5_SIG, ROM11_DATA6_SIG, ROM11_DATA7_SIG, ROM11_DATA8_SIG, ROM11_DATA9_SIG,
       ROM11_DATA10_SIG, ROM11_DATA11_SIG, ROM11_DATA12_SIG, ROM11_DATA13_SIG, ROM11_DATA14_SIG,
       ROM11_DATA15_SIG, ROM11_DATA16_SIG, ROM11_DATA17_SIG, ROM11_DATA18_SIG, ROM11_DATA19_SIG,
       ROM11_DATA20_SIG, ROM11_DATA21_SIG, ROM11_DATA22_SIG, ROM11_DATA23_SIG, ROM11_DATA24_SIG, ROM11_DATA25_SIG,
       ROM11_DATA26_SIG, ROM11_DATA27_SIG, ROM11_DATA28_SIG, ROM11_DATA29_SIG, ROM11_DATA30_SIG, ROM11_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM12_DATA0_SIG, ROM12_DATA1_SIG, ROM12_DATA2_SIG, ROM12_DATA3_SIG, ROM12_DATA4_SIG,
       ROM12_DATA5_SIG, ROM12_DATA6_SIG, ROM12_DATA7_SIG, ROM12_DATA8_SIG, ROM12_DATA9_SIG,
       ROM12_DATA10_SIG, ROM12_DATA11_SIG, ROM12_DATA12_SIG, ROM12_DATA13_SIG, ROM12_DATA14_SIG,
       ROM12_DATA15_SIG, ROM12_DATA16_SIG, ROM12_DATA17_SIG, ROM12_DATA18_SIG, ROM12_DATA19_SIG,
       ROM12_DATA20_SIG, ROM12_DATA21_SIG, ROM12_DATA22_SIG, ROM12_DATA23_SIG, ROM12_DATA24_SIG, ROM12_DATA25_SIG,
       ROM12_DATA26_SIG, ROM12_DATA27_SIG, ROM12_DATA28_SIG, ROM12_DATA29_SIG, ROM12_DATA30_SIG, ROM12_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM13_DATA0_SIG, ROM13_DATA1_SIG, ROM13_DATA2_SIG, ROM13_DATA3_SIG, ROM13_DATA4_SIG,
       ROM13_DATA5_SIG, ROM13_DATA6_SIG, ROM13_DATA7_SIG, ROM13_DATA8_SIG, ROM13_DATA9_SIG,
       ROM13_DATA10_SIG, ROM13_DATA11_SIG, ROM13_DATA12_SIG, ROM13_DATA13_SIG, ROM13_DATA14_SIG,
       ROM13_DATA15_SIG, ROM13_DATA16_SIG, ROM13_DATA17_SIG, ROM13_DATA18_SIG, ROM13_DATA19_SIG,
       ROM13_DATA20_SIG, ROM13_DATA21_SIG, ROM13_DATA22_SIG, ROM13_DATA23_SIG, ROM13_DATA24_SIG, ROM13_DATA25_SIG,
       ROM13_DATA26_SIG, ROM13_DATA27_SIG, ROM13_DATA28_SIG, ROM13_DATA29_SIG, ROM13_DATA30_SIG, ROM13_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM14_DATA0_SIG, ROM14_DATA1_SIG, ROM14_DATA2_SIG, ROM14_DATA3_SIG, ROM14_DATA4_SIG,
       ROM14_DATA5_SIG, ROM14_DATA6_SIG, ROM14_DATA7_SIG, ROM14_DATA8_SIG, ROM14_DATA9_SIG,
       ROM14_DATA10_SIG, ROM14_DATA11_SIG, ROM14_DATA12_SIG, ROM14_DATA13_SIG, ROM14_DATA14_SIG,
       ROM14_DATA15_SIG, ROM14_DATA16_SIG, ROM14_DATA17_SIG, ROM14_DATA18_SIG, ROM14_DATA19_SIG,
       ROM14_DATA20_SIG, ROM14_DATA21_SIG, ROM14_DATA22_SIG, ROM14_DATA23_SIG, ROM14_DATA24_SIG, ROM14_DATA25_SIG,
       ROM14_DATA26_SIG, ROM14_DATA27_SIG, ROM14_DATA28_SIG, ROM14_DATA29_SIG, ROM14_DATA30_SIG, ROM14_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM15_DATA0_SIG, ROM15_DATA1_SIG, ROM15_DATA2_SIG, ROM15_DATA3_SIG, ROM15_DATA4_SIG,
       ROM15_DATA5_SIG, ROM15_DATA6_SIG, ROM15_DATA7_SIG, ROM15_DATA8_SIG, ROM15_DATA9_SIG,
       ROM15_DATA10_SIG, ROM15_DATA11_SIG, ROM15_DATA12_SIG, ROM15_DATA13_SIG, ROM15_DATA14_SIG,
       ROM15_DATA15_SIG, ROM15_DATA16_SIG, ROM15_DATA17_SIG, ROM15_DATA18_SIG, ROM15_DATA19_SIG,
       ROM15_DATA20_SIG, ROM15_DATA21_SIG, ROM15_DATA22_SIG, ROM15_DATA23_SIG, ROM15_DATA24_SIG, ROM15_DATA25_SIG,
       ROM15_DATA26_SIG, ROM15_DATA27_SIG, ROM15_DATA28_SIG, ROM15_DATA29_SIG, ROM15_DATA30_SIG, ROM15_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM16_DATA0_SIG, ROM16_DATA1_SIG, ROM16_DATA2_SIG, ROM16_DATA3_SIG, ROM16_DATA4_SIG,
       ROM16_DATA5_SIG, ROM16_DATA6_SIG, ROM16_DATA7_SIG, ROM16_DATA8_SIG, ROM16_DATA9_SIG,
       ROM16_DATA10_SIG, ROM16_DATA11_SIG, ROM16_DATA12_SIG, ROM16_DATA13_SIG, ROM16_DATA14_SIG,
       ROM16_DATA15_SIG, ROM16_DATA16_SIG, ROM16_DATA17_SIG, ROM16_DATA18_SIG, ROM16_DATA19_SIG,
       ROM16_DATA20_SIG, ROM16_DATA21_SIG, ROM16_DATA22_SIG, ROM16_DATA23_SIG, ROM16_DATA24_SIG, ROM16_DATA25_SIG,
       ROM16_DATA26_SIG, ROM16_DATA27_SIG, ROM16_DATA28_SIG, ROM16_DATA29_SIG, ROM16_DATA30_SIG, ROM16_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM17_DATA0_SIG, ROM17_DATA1_SIG, ROM17_DATA2_SIG, ROM17_DATA3_SIG, ROM17_DATA4_SIG,
       ROM17_DATA5_SIG, ROM17_DATA6_SIG, ROM17_DATA7_SIG, ROM17_DATA8_SIG, ROM17_DATA9_SIG,
       ROM17_DATA10_SIG, ROM17_DATA11_SIG, ROM17_DATA12_SIG, ROM17_DATA13_SIG, ROM17_DATA14_SIG,
       ROM17_DATA15_SIG, ROM17_DATA16_SIG, ROM17_DATA17_SIG, ROM17_DATA18_SIG, ROM17_DATA19_SIG,
       ROM17_DATA20_SIG, ROM17_DATA21_SIG, ROM17_DATA22_SIG, ROM17_DATA23_SIG, ROM17_DATA24_SIG, ROM17_DATA25_SIG,
       ROM17_DATA26_SIG, ROM17_DATA27_SIG, ROM17_DATA28_SIG, ROM17_DATA29_SIG, ROM17_DATA30_SIG, ROM17_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM18_DATA0_SIG, ROM18_DATA1_SIG, ROM18_DATA2_SIG, ROM18_DATA3_SIG, ROM18_DATA4_SIG,
       ROM18_DATA5_SIG, ROM18_DATA6_SIG, ROM18_DATA7_SIG, ROM18_DATA8_SIG, ROM18_DATA9_SIG,
       ROM18_DATA10_SIG, ROM18_DATA11_SIG, ROM18_DATA12_SIG, ROM18_DATA13_SIG, ROM18_DATA14_SIG,
       ROM18_DATA15_SIG, ROM18_DATA16_SIG, ROM18_DATA17_SIG, ROM18_DATA18_SIG, ROM18_DATA19_SIG,
       ROM18_DATA20_SIG, ROM18_DATA21_SIG, ROM18_DATA22_SIG, ROM18_DATA23_SIG, ROM18_DATA24_SIG, ROM18_DATA25_SIG,
       ROM18_DATA26_SIG, ROM18_DATA27_SIG, ROM18_DATA28_SIG, ROM18_DATA29_SIG, ROM18_DATA30_SIG, ROM18_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM19_DATA0_SIG, ROM19_DATA1_SIG, ROM19_DATA2_SIG, ROM19_DATA3_SIG, ROM19_DATA4_SIG,
       ROM19_DATA5_SIG, ROM19_DATA6_SIG, ROM19_DATA7_SIG, ROM19_DATA8_SIG, ROM19_DATA9_SIG,
       ROM19_DATA10_SIG, ROM19_DATA11_SIG, ROM19_DATA12_SIG, ROM19_DATA13_SIG, ROM19_DATA14_SIG,
       ROM19_DATA15_SIG, ROM19_DATA16_SIG, ROM19_DATA17_SIG, ROM19_DATA18_SIG, ROM19_DATA19_SIG,
       ROM19_DATA20_SIG, ROM19_DATA21_SIG, ROM19_DATA22_SIG, ROM19_DATA23_SIG, ROM19_DATA24_SIG, ROM19_DATA25_SIG,
       ROM19_DATA26_SIG, ROM19_DATA27_SIG, ROM19_DATA28_SIG, ROM19_DATA29_SIG, ROM19_DATA30_SIG, ROM19_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM20_DATA0_SIG, ROM20_DATA1_SIG, ROM20_DATA2_SIG, ROM20_DATA3_SIG, ROM20_DATA4_SIG,
       ROM20_DATA5_SIG, ROM20_DATA6_SIG, ROM20_DATA7_SIG, ROM20_DATA8_SIG, ROM20_DATA9_SIG,
       ROM20_DATA10_SIG, ROM20_DATA11_SIG, ROM20_DATA12_SIG, ROM20_DATA13_SIG, ROM20_DATA14_SIG,
       ROM20_DATA15_SIG, ROM20_DATA16_SIG, ROM20_DATA17_SIG, ROM20_DATA18_SIG, ROM20_DATA19_SIG,
       ROM20_DATA20_SIG, ROM20_DATA21_SIG, ROM20_DATA22_SIG, ROM20_DATA23_SIG, ROM20_DATA24_SIG, ROM20_DATA25_SIG,
       ROM20_DATA26_SIG, ROM20_DATA27_SIG, ROM20_DATA28_SIG, ROM20_DATA29_SIG, ROM20_DATA30_SIG, ROM20_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM21_DATA0_SIG, ROM21_DATA1_SIG, ROM21_DATA2_SIG, ROM21_DATA3_SIG, ROM21_DATA4_SIG,
       ROM21_DATA5_SIG, ROM21_DATA6_SIG, ROM21_DATA7_SIG, ROM21_DATA8_SIG, ROM21_DATA9_SIG,
       ROM21_DATA10_SIG, ROM21_DATA11_SIG, ROM21_DATA12_SIG, ROM21_DATA13_SIG, ROM21_DATA14_SIG,
       ROM21_DATA15_SIG, ROM21_DATA16_SIG, ROM21_DATA17_SIG, ROM21_DATA18_SIG, ROM21_DATA19_SIG,
       ROM21_DATA20_SIG, ROM21_DATA21_SIG, ROM21_DATA22_SIG, ROM21_DATA23_SIG, ROM21_DATA24_SIG, ROM21_DATA25_SIG,
       ROM21_DATA26_SIG, ROM21_DATA27_SIG, ROM21_DATA28_SIG, ROM21_DATA29_SIG, ROM21_DATA30_SIG, ROM21_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM22_DATA0_SIG, ROM22_DATA1_SIG, ROM22_DATA2_SIG, ROM22_DATA3_SIG, ROM22_DATA4_SIG,
       ROM22_DATA5_SIG, ROM22_DATA6_SIG, ROM22_DATA7_SIG, ROM22_DATA8_SIG, ROM22_DATA9_SIG,
       ROM22_DATA10_SIG, ROM22_DATA11_SIG, ROM22_DATA12_SIG, ROM22_DATA13_SIG, ROM22_DATA14_SIG,
       ROM22_DATA15_SIG, ROM22_DATA16_SIG, ROM22_DATA17_SIG, ROM22_DATA18_SIG, ROM22_DATA19_SIG,
       ROM22_DATA20_SIG, ROM22_DATA21_SIG, ROM22_DATA22_SIG, ROM22_DATA23_SIG, ROM22_DATA24_SIG, ROM22_DATA25_SIG,
       ROM22_DATA26_SIG, ROM22_DATA27_SIG, ROM22_DATA28_SIG, ROM22_DATA29_SIG, ROM22_DATA30_SIG, ROM22_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM23_DATA0_SIG, ROM23_DATA1_SIG, ROM23_DATA2_SIG, ROM23_DATA3_SIG, ROM23_DATA4_SIG,
       ROM23_DATA5_SIG, ROM23_DATA6_SIG, ROM23_DATA7_SIG, ROM23_DATA8_SIG, ROM23_DATA9_SIG,
       ROM23_DATA10_SIG, ROM23_DATA11_SIG, ROM23_DATA12_SIG, ROM23_DATA13_SIG, ROM23_DATA14_SIG,
       ROM23_DATA15_SIG, ROM23_DATA16_SIG, ROM23_DATA17_SIG, ROM23_DATA18_SIG, ROM23_DATA19_SIG,
       ROM23_DATA20_SIG, ROM23_DATA21_SIG, ROM23_DATA22_SIG, ROM23_DATA23_SIG, ROM23_DATA24_SIG, ROM23_DATA25_SIG,
       ROM23_DATA26_SIG, ROM23_DATA27_SIG, ROM23_DATA28_SIG, ROM23_DATA29_SIG, ROM23_DATA30_SIG, ROM23_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM24_DATA0_SIG, ROM24_DATA1_SIG, ROM24_DATA2_SIG, ROM24_DATA3_SIG, ROM24_DATA4_SIG,
       ROM24_DATA5_SIG, ROM24_DATA6_SIG, ROM24_DATA7_SIG, ROM24_DATA8_SIG, ROM24_DATA9_SIG,
       ROM24_DATA10_SIG, ROM24_DATA11_SIG, ROM24_DATA12_SIG, ROM24_DATA13_SIG, ROM24_DATA14_SIG,
       ROM24_DATA15_SIG, ROM24_DATA16_SIG, ROM24_DATA17_SIG, ROM24_DATA18_SIG, ROM24_DATA19_SIG,
       ROM24_DATA20_SIG, ROM24_DATA21_SIG, ROM24_DATA22_SIG, ROM24_DATA23_SIG, ROM24_DATA24_SIG, ROM24_DATA25_SIG,
       ROM24_DATA26_SIG, ROM24_DATA27_SIG, ROM24_DATA28_SIG, ROM24_DATA29_SIG, ROM24_DATA30_SIG, ROM24_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM25_DATA0_SIG, ROM25_DATA1_SIG, ROM25_DATA2_SIG, ROM25_DATA3_SIG, ROM25_DATA4_SIG,
       ROM25_DATA5_SIG, ROM25_DATA6_SIG, ROM25_DATA7_SIG, ROM25_DATA8_SIG, ROM25_DATA9_SIG,
       ROM25_DATA10_SIG, ROM25_DATA11_SIG, ROM25_DATA12_SIG, ROM25_DATA13_SIG, ROM25_DATA14_SIG,
       ROM25_DATA15_SIG, ROM25_DATA16_SIG, ROM25_DATA17_SIG, ROM25_DATA18_SIG, ROM25_DATA19_SIG,
       ROM25_DATA20_SIG, ROM25_DATA21_SIG, ROM25_DATA22_SIG, ROM25_DATA23_SIG, ROM25_DATA24_SIG, ROM25_DATA25_SIG,
       ROM25_DATA26_SIG, ROM25_DATA27_SIG, ROM25_DATA28_SIG, ROM25_DATA29_SIG, ROM25_DATA30_SIG, ROM25_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM26_DATA0_SIG, ROM26_DATA1_SIG, ROM26_DATA2_SIG, ROM26_DATA3_SIG, ROM26_DATA4_SIG,
       ROM26_DATA5_SIG, ROM26_DATA6_SIG, ROM26_DATA7_SIG, ROM26_DATA8_SIG, ROM26_DATA9_SIG,
       ROM26_DATA10_SIG, ROM26_DATA11_SIG, ROM26_DATA12_SIG, ROM26_DATA13_SIG, ROM26_DATA14_SIG,
       ROM26_DATA15_SIG, ROM26_DATA16_SIG, ROM26_DATA17_SIG, ROM26_DATA18_SIG, ROM26_DATA19_SIG,
       ROM26_DATA20_SIG, ROM26_DATA21_SIG, ROM26_DATA22_SIG, ROM26_DATA23_SIG, ROM26_DATA24_SIG, ROM26_DATA25_SIG,
       ROM26_DATA26_SIG, ROM26_DATA27_SIG, ROM26_DATA28_SIG, ROM26_DATA29_SIG, ROM26_DATA30_SIG, ROM26_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM27_DATA0_SIG, ROM27_DATA1_SIG, ROM27_DATA2_SIG, ROM27_DATA3_SIG, ROM27_DATA4_SIG,
       ROM27_DATA5_SIG, ROM27_DATA6_SIG, ROM27_DATA7_SIG, ROM27_DATA8_SIG, ROM27_DATA9_SIG,
       ROM27_DATA10_SIG, ROM27_DATA11_SIG, ROM27_DATA12_SIG, ROM27_DATA13_SIG, ROM27_DATA14_SIG,
       ROM27_DATA15_SIG, ROM27_DATA16_SIG, ROM27_DATA17_SIG, ROM27_DATA18_SIG, ROM27_DATA19_SIG,
       ROM27_DATA20_SIG, ROM27_DATA21_SIG, ROM27_DATA22_SIG, ROM27_DATA23_SIG, ROM27_DATA24_SIG, ROM27_DATA25_SIG,
       ROM27_DATA26_SIG, ROM27_DATA27_SIG, ROM27_DATA28_SIG, ROM27_DATA29_SIG, ROM27_DATA30_SIG, ROM27_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM28_DATA0_SIG, ROM28_DATA1_SIG, ROM28_DATA2_SIG, ROM28_DATA3_SIG, ROM28_DATA4_SIG,
       ROM28_DATA5_SIG, ROM28_DATA6_SIG, ROM28_DATA7_SIG, ROM28_DATA8_SIG, ROM28_DATA9_SIG,
       ROM28_DATA10_SIG, ROM28_DATA11_SIG, ROM28_DATA12_SIG, ROM28_DATA13_SIG, ROM28_DATA14_SIG,
       ROM28_DATA15_SIG, ROM28_DATA16_SIG, ROM28_DATA17_SIG, ROM28_DATA18_SIG, ROM28_DATA19_SIG,
       ROM28_DATA20_SIG, ROM28_DATA21_SIG, ROM28_DATA22_SIG, ROM28_DATA23_SIG, ROM28_DATA24_SIG, ROM28_DATA25_SIG,
       ROM28_DATA26_SIG, ROM28_DATA27_SIG, ROM28_DATA28_SIG, ROM28_DATA29_SIG, ROM28_DATA30_SIG, ROM28_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM29_DATA0_SIG, ROM29_DATA1_SIG, ROM29_DATA2_SIG, ROM29_DATA3_SIG, ROM29_DATA4_SIG,
       ROM29_DATA5_SIG, ROM29_DATA6_SIG, ROM29_DATA7_SIG, ROM29_DATA8_SIG, ROM29_DATA9_SIG,
       ROM29_DATA10_SIG, ROM29_DATA11_SIG, ROM29_DATA12_SIG, ROM29_DATA13_SIG, ROM29_DATA14_SIG,
       ROM29_DATA15_SIG, ROM29_DATA16_SIG, ROM29_DATA17_SIG, ROM29_DATA18_SIG, ROM29_DATA19_SIG,
       ROM29_DATA20_SIG, ROM29_DATA21_SIG, ROM29_DATA22_SIG, ROM29_DATA23_SIG, ROM29_DATA24_SIG, ROM29_DATA25_SIG,
       ROM29_DATA26_SIG, ROM29_DATA27_SIG, ROM29_DATA28_SIG, ROM29_DATA29_SIG, ROM29_DATA30_SIG, ROM29_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM30_DATA0_SIG, ROM30_DATA1_SIG, ROM30_DATA2_SIG, ROM30_DATA3_SIG, ROM30_DATA4_SIG,
       ROM30_DATA5_SIG, ROM30_DATA6_SIG, ROM30_DATA7_SIG, ROM30_DATA8_SIG, ROM30_DATA9_SIG,
       ROM30_DATA10_SIG, ROM30_DATA11_SIG, ROM30_DATA12_SIG, ROM30_DATA13_SIG, ROM30_DATA14_SIG,
       ROM30_DATA15_SIG, ROM30_DATA16_SIG, ROM30_DATA17_SIG, ROM30_DATA18_SIG, ROM30_DATA19_SIG,
       ROM30_DATA20_SIG, ROM30_DATA21_SIG, ROM30_DATA22_SIG, ROM30_DATA23_SIG, ROM30_DATA24_SIG, ROM30_DATA25_SIG,
       ROM30_DATA26_SIG, ROM30_DATA27_SIG, ROM30_DATA28_SIG, ROM30_DATA29_SIG, ROM30_DATA30_SIG, ROM30_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM31_DATA0_SIG, ROM31_DATA1_SIG, ROM31_DATA2_SIG, ROM31_DATA3_SIG, ROM31_DATA4_SIG,
       ROM31_DATA5_SIG, ROM31_DATA6_SIG, ROM31_DATA7_SIG, ROM31_DATA8_SIG, ROM31_DATA9_SIG,
       ROM31_DATA10_SIG, ROM31_DATA11_SIG, ROM31_DATA12_SIG, ROM31_DATA13_SIG, ROM31_DATA14_SIG,
       ROM31_DATA15_SIG, ROM31_DATA16_SIG, ROM31_DATA17_SIG, ROM31_DATA18_SIG, ROM31_DATA19_SIG,
       ROM31_DATA20_SIG, ROM31_DATA21_SIG, ROM31_DATA22_SIG, ROM31_DATA23_SIG, ROM31_DATA24_SIG, ROM31_DATA25_SIG,
       ROM31_DATA26_SIG, ROM31_DATA27_SIG, ROM31_DATA28_SIG, ROM31_DATA29_SIG, ROM31_DATA30_SIG, ROM31_DATA31_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');

signal ADDR0_0_SIG, ADDR0_1_SIG, ADDR0_2_SIG, ADDR0_3_SIG, ADDR0_4_SIG, ADDR0_5_SIG, ADDR0_6_SIG, ADDR0_7_SIG,
       ADDR0_8_SIG, ADDR0_9_SIG, ADDR0_10_SIG, ADDR0_11_SIG, ADDR0_12_SIG, ADDR0_13_SIG, ADDR0_14_SIG, ADDR0_15_SIG,
       ADDR0_16_SIG, ADDR0_17_SIG, ADDR0_18_SIG, ADDR0_19_SIG, ADDR0_20_SIG, ADDR0_21_SIG, ADDR0_22_SIG, ADDR0_23_SIG,
       ADDR0_24_SIG, ADDR0_25_SIG, ADDR0_26_SIG, ADDR0_27_SIG, ADDR0_28_SIG, ADDR0_29_SIG, ADDR0_30_SIG, ADDR0_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR1_0_SIG, ADDR1_1_SIG, ADDR1_2_SIG, ADDR1_3_SIG, ADDR1_4_SIG, ADDR1_5_SIG, ADDR1_6_SIG, ADDR1_7_SIG,
       ADDR1_8_SIG, ADDR1_9_SIG, ADDR1_10_SIG, ADDR1_11_SIG, ADDR1_12_SIG, ADDR1_13_SIG, ADDR1_14_SIG, ADDR1_15_SIG,
       ADDR1_16_SIG, ADDR1_17_SIG, ADDR1_18_SIG, ADDR1_19_SIG, ADDR1_20_SIG, ADDR1_21_SIG, ADDR1_22_SIG, ADDR1_23_SIG,
       ADDR1_24_SIG, ADDR1_25_SIG, ADDR1_26_SIG, ADDR1_27_SIG, ADDR1_28_SIG, ADDR1_29_SIG, ADDR1_30_SIG, ADDR1_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR2_0_SIG, ADDR2_1_SIG, ADDR2_2_SIG, ADDR2_3_SIG, ADDR2_4_SIG, ADDR2_5_SIG, ADDR2_6_SIG, ADDR2_7_SIG,
       ADDR2_8_SIG, ADDR2_9_SIG, ADDR2_10_SIG, ADDR2_11_SIG, ADDR2_12_SIG, ADDR2_13_SIG, ADDR2_14_SIG, ADDR2_15_SIG,
       ADDR2_16_SIG, ADDR2_17_SIG, ADDR2_18_SIG, ADDR2_19_SIG, ADDR2_20_SIG, ADDR2_21_SIG, ADDR2_22_SIG, ADDR2_23_SIG,
       ADDR2_24_SIG, ADDR2_25_SIG, ADDR2_26_SIG, ADDR2_27_SIG, ADDR2_28_SIG, ADDR2_29_SIG, ADDR2_30_SIG, ADDR2_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR3_0_SIG, ADDR3_1_SIG, ADDR3_2_SIG, ADDR3_3_SIG, ADDR3_4_SIG, ADDR3_5_SIG, ADDR3_6_SIG, ADDR3_7_SIG,
       ADDR3_8_SIG, ADDR3_9_SIG, ADDR3_10_SIG, ADDR3_11_SIG, ADDR3_12_SIG, ADDR3_13_SIG, ADDR3_14_SIG, ADDR3_15_SIG,
       ADDR3_16_SIG, ADDR3_17_SIG, ADDR3_18_SIG, ADDR3_19_SIG, ADDR3_20_SIG, ADDR3_21_SIG, ADDR3_22_SIG, ADDR3_23_SIG,
       ADDR3_24_SIG, ADDR3_25_SIG, ADDR3_26_SIG, ADDR3_27_SIG, ADDR3_28_SIG, ADDR3_29_SIG, ADDR3_30_SIG, ADDR3_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR4_0_SIG, ADDR4_1_SIG, ADDR4_2_SIG, ADDR4_3_SIG, ADDR4_4_SIG, ADDR4_5_SIG, ADDR4_6_SIG, ADDR4_7_SIG,
       ADDR4_8_SIG, ADDR4_9_SIG, ADDR4_10_SIG, ADDR4_11_SIG, ADDR4_12_SIG, ADDR4_13_SIG, ADDR4_14_SIG, ADDR4_15_SIG,
       ADDR4_16_SIG, ADDR4_17_SIG, ADDR4_18_SIG, ADDR4_19_SIG, ADDR4_20_SIG, ADDR4_21_SIG, ADDR4_22_SIG, ADDR4_23_SIG,
       ADDR4_24_SIG, ADDR4_25_SIG, ADDR4_26_SIG, ADDR4_27_SIG, ADDR4_28_SIG, ADDR4_29_SIG, ADDR4_30_SIG, ADDR4_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR5_0_SIG, ADDR5_1_SIG, ADDR5_2_SIG, ADDR5_3_SIG, ADDR5_4_SIG, ADDR5_5_SIG, ADDR5_6_SIG, ADDR5_7_SIG,
       ADDR5_8_SIG, ADDR5_9_SIG, ADDR5_10_SIG, ADDR5_11_SIG, ADDR5_12_SIG, ADDR5_13_SIG, ADDR5_14_SIG, ADDR5_15_SIG,
       ADDR5_16_SIG, ADDR5_17_SIG, ADDR5_18_SIG, ADDR5_19_SIG, ADDR5_20_SIG, ADDR5_21_SIG, ADDR5_22_SIG, ADDR5_23_SIG,
       ADDR5_24_SIG, ADDR5_25_SIG, ADDR5_26_SIG, ADDR5_27_SIG, ADDR5_28_SIG, ADDR5_29_SIG, ADDR5_30_SIG, ADDR5_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR6_0_SIG, ADDR6_1_SIG, ADDR6_2_SIG, ADDR6_3_SIG, ADDR6_4_SIG, ADDR6_5_SIG, ADDR6_6_SIG, ADDR6_7_SIG,
       ADDR6_8_SIG, ADDR6_9_SIG, ADDR6_10_SIG, ADDR6_11_SIG, ADDR6_12_SIG, ADDR6_13_SIG, ADDR6_14_SIG, ADDR6_15_SIG,
       ADDR6_16_SIG, ADDR6_17_SIG, ADDR6_18_SIG, ADDR6_19_SIG, ADDR6_20_SIG, ADDR6_21_SIG, ADDR6_22_SIG, ADDR6_23_SIG,
       ADDR6_24_SIG, ADDR6_25_SIG, ADDR6_26_SIG, ADDR6_27_SIG, ADDR6_28_SIG, ADDR6_29_SIG, ADDR6_30_SIG, ADDR6_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR7_0_SIG, ADDR7_1_SIG, ADDR7_2_SIG, ADDR7_3_SIG, ADDR7_4_SIG, ADDR7_5_SIG, ADDR7_6_SIG, ADDR7_7_SIG,
       ADDR7_8_SIG, ADDR7_9_SIG, ADDR7_10_SIG, ADDR7_11_SIG, ADDR7_12_SIG, ADDR7_13_SIG, ADDR7_14_SIG, ADDR7_15_SIG,
       ADDR7_16_SIG, ADDR7_17_SIG, ADDR7_18_SIG, ADDR7_19_SIG, ADDR7_20_SIG, ADDR7_21_SIG, ADDR7_22_SIG, ADDR7_23_SIG,
       ADDR7_24_SIG, ADDR7_25_SIG, ADDR7_26_SIG, ADDR7_27_SIG, ADDR7_28_SIG, ADDR7_29_SIG, ADDR7_30_SIG, ADDR7_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR8_0_SIG, ADDR8_1_SIG, ADDR8_2_SIG, ADDR8_3_SIG, ADDR8_4_SIG, ADDR8_5_SIG, ADDR8_6_SIG, ADDR8_7_SIG,
       ADDR8_8_SIG, ADDR8_9_SIG, ADDR8_10_SIG, ADDR8_11_SIG, ADDR8_12_SIG, ADDR8_13_SIG, ADDR8_14_SIG, ADDR8_15_SIG,
       ADDR8_16_SIG, ADDR8_17_SIG, ADDR8_18_SIG, ADDR8_19_SIG, ADDR8_20_SIG, ADDR8_21_SIG, ADDR8_22_SIG, ADDR8_23_SIG,
       ADDR8_24_SIG, ADDR8_25_SIG, ADDR8_26_SIG, ADDR8_27_SIG, ADDR8_28_SIG, ADDR8_29_SIG, ADDR8_30_SIG, ADDR8_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR9_0_SIG, ADDR9_1_SIG, ADDR9_2_SIG, ADDR9_3_SIG, ADDR9_4_SIG, ADDR9_5_SIG, ADDR9_6_SIG, ADDR9_7_SIG,
       ADDR9_8_SIG, ADDR9_9_SIG, ADDR9_10_SIG, ADDR9_11_SIG, ADDR9_12_SIG, ADDR9_13_SIG, ADDR9_14_SIG, ADDR9_15_SIG,
       ADDR9_16_SIG, ADDR9_17_SIG, ADDR9_18_SIG, ADDR9_19_SIG, ADDR9_20_SIG, ADDR9_21_SIG, ADDR9_22_SIG, ADDR9_23_SIG,
       ADDR9_24_SIG, ADDR9_25_SIG, ADDR9_26_SIG, ADDR9_27_SIG, ADDR9_28_SIG, ADDR9_29_SIG, ADDR9_30_SIG, ADDR9_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR10_0_SIG, ADDR10_1_SIG, ADDR10_2_SIG, ADDR10_3_SIG, ADDR10_4_SIG, ADDR10_5_SIG, ADDR10_6_SIG, ADDR10_7_SIG,
       ADDR10_8_SIG, ADDR10_9_SIG, ADDR10_10_SIG, ADDR10_11_SIG, ADDR10_12_SIG, ADDR10_13_SIG, ADDR10_14_SIG, ADDR10_15_SIG,
       ADDR10_16_SIG, ADDR10_17_SIG, ADDR10_18_SIG, ADDR10_19_SIG, ADDR10_20_SIG, ADDR10_21_SIG, ADDR10_22_SIG, ADDR10_23_SIG,
       ADDR10_24_SIG, ADDR10_25_SIG, ADDR10_26_SIG, ADDR10_27_SIG, ADDR10_28_SIG, ADDR10_29_SIG, ADDR10_30_SIG, ADDR10_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR11_0_SIG, ADDR11_1_SIG, ADDR11_2_SIG, ADDR11_3_SIG, ADDR11_4_SIG, ADDR11_5_SIG, ADDR11_6_SIG, ADDR11_7_SIG,
       ADDR11_8_SIG, ADDR11_9_SIG, ADDR11_10_SIG, ADDR11_11_SIG, ADDR11_12_SIG, ADDR11_13_SIG, ADDR11_14_SIG, ADDR11_15_SIG,
       ADDR11_16_SIG, ADDR11_17_SIG, ADDR11_18_SIG, ADDR11_19_SIG, ADDR11_20_SIG, ADDR11_21_SIG, ADDR11_22_SIG, ADDR11_23_SIG,
       ADDR11_24_SIG, ADDR11_25_SIG, ADDR11_26_SIG, ADDR11_27_SIG, ADDR11_28_SIG, ADDR11_29_SIG, ADDR11_30_SIG, ADDR11_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR12_0_SIG, ADDR12_1_SIG, ADDR12_2_SIG, ADDR12_3_SIG, ADDR12_4_SIG, ADDR12_5_SIG, ADDR12_6_SIG, ADDR12_7_SIG,
       ADDR12_8_SIG, ADDR12_9_SIG, ADDR12_10_SIG, ADDR12_11_SIG, ADDR12_12_SIG, ADDR12_13_SIG, ADDR12_14_SIG, ADDR12_15_SIG,
       ADDR12_16_SIG, ADDR12_17_SIG, ADDR12_18_SIG, ADDR12_19_SIG, ADDR12_20_SIG, ADDR12_21_SIG, ADDR12_22_SIG, ADDR12_23_SIG,
       ADDR12_24_SIG, ADDR12_25_SIG, ADDR12_26_SIG, ADDR12_27_SIG, ADDR12_28_SIG, ADDR12_29_SIG, ADDR12_30_SIG, ADDR12_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR13_0_SIG, ADDR13_1_SIG, ADDR13_2_SIG, ADDR13_3_SIG, ADDR13_4_SIG, ADDR13_5_SIG, ADDR13_6_SIG, ADDR13_7_SIG,
       ADDR13_8_SIG, ADDR13_9_SIG, ADDR13_10_SIG, ADDR13_11_SIG, ADDR13_12_SIG, ADDR13_13_SIG, ADDR13_14_SIG, ADDR13_15_SIG,
       ADDR13_16_SIG, ADDR13_17_SIG, ADDR13_18_SIG, ADDR13_19_SIG, ADDR13_20_SIG, ADDR13_21_SIG, ADDR13_22_SIG, ADDR13_23_SIG,
       ADDR13_24_SIG, ADDR13_25_SIG, ADDR13_26_SIG, ADDR13_27_SIG, ADDR13_28_SIG, ADDR13_29_SIG, ADDR13_30_SIG, ADDR13_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR14_0_SIG, ADDR14_1_SIG, ADDR14_2_SIG, ADDR14_3_SIG, ADDR14_4_SIG, ADDR14_5_SIG, ADDR14_6_SIG, ADDR14_7_SIG,
       ADDR14_8_SIG, ADDR14_9_SIG, ADDR14_10_SIG, ADDR14_11_SIG, ADDR14_12_SIG, ADDR14_13_SIG, ADDR14_14_SIG, ADDR14_15_SIG,
       ADDR14_16_SIG, ADDR14_17_SIG, ADDR14_18_SIG, ADDR14_19_SIG, ADDR14_20_SIG, ADDR14_21_SIG, ADDR14_22_SIG, ADDR14_23_SIG,
       ADDR14_24_SIG, ADDR14_25_SIG, ADDR14_26_SIG, ADDR14_27_SIG, ADDR14_28_SIG, ADDR14_29_SIG, ADDR14_30_SIG, ADDR14_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR15_0_SIG, ADDR15_1_SIG, ADDR15_2_SIG, ADDR15_3_SIG, ADDR15_4_SIG, ADDR15_5_SIG, ADDR15_6_SIG, ADDR15_7_SIG,
       ADDR15_8_SIG, ADDR15_9_SIG, ADDR15_10_SIG, ADDR15_11_SIG, ADDR15_12_SIG, ADDR15_13_SIG, ADDR15_14_SIG, ADDR15_15_SIG,
       ADDR15_16_SIG, ADDR15_17_SIG, ADDR15_18_SIG, ADDR15_19_SIG, ADDR15_20_SIG, ADDR15_21_SIG, ADDR15_22_SIG, ADDR15_23_SIG,
       ADDR15_24_SIG, ADDR15_25_SIG, ADDR15_26_SIG, ADDR15_27_SIG, ADDR15_28_SIG, ADDR15_29_SIG, ADDR15_30_SIG, ADDR15_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR16_0_SIG, ADDR16_1_SIG, ADDR16_2_SIG,  ADDR16_3_SIG,  ADDR16_4_SIG,  ADDR16_5_SIG,  ADDR16_6_SIG,  ADDR16_7_SIG,
       ADDR16_8_SIG, ADDR16_9_SIG, ADDR16_10_SIG, ADDR16_11_SIG, ADDR16_12_SIG, ADDR16_13_SIG, ADDR16_14_SIG, ADDR16_15_SIG,
       ADDR16_16_SIG, ADDR16_17_SIG, ADDR16_18_SIG, ADDR16_19_SIG, ADDR16_20_SIG, ADDR16_21_SIG, ADDR16_22_SIG, ADDR16_23_SIG,
       ADDR16_24_SIG, ADDR16_25_SIG, ADDR16_26_SIG, ADDR16_27_SIG, ADDR16_28_SIG, ADDR16_29_SIG, ADDR16_30_SIG, ADDR16_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR17_0_SIG, ADDR17_1_SIG, ADDR17_2_SIG,  ADDR17_3_SIG,  ADDR17_4_SIG,  ADDR17_5_SIG,  ADDR17_6_SIG,  ADDR17_7_SIG,
       ADDR17_8_SIG, ADDR17_9_SIG, ADDR17_10_SIG, ADDR17_11_SIG, ADDR17_12_SIG, ADDR17_13_SIG, ADDR17_14_SIG, ADDR17_15_SIG,
       ADDR17_16_SIG, ADDR17_17_SIG, ADDR17_18_SIG, ADDR17_19_SIG, ADDR17_20_SIG, ADDR17_21_SIG, ADDR17_22_SIG, ADDR17_23_SIG,
       ADDR17_24_SIG, ADDR17_25_SIG, ADDR17_26_SIG, ADDR17_27_SIG, ADDR17_28_SIG, ADDR17_29_SIG, ADDR17_30_SIG, ADDR17_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR18_0_SIG, ADDR18_1_SIG, ADDR18_2_SIG,  ADDR18_3_SIG,  ADDR18_4_SIG,  ADDR18_5_SIG,  ADDR18_6_SIG,  ADDR18_7_SIG,
       ADDR18_8_SIG, ADDR18_9_SIG, ADDR18_10_SIG, ADDR18_11_SIG, ADDR18_12_SIG, ADDR18_13_SIG, ADDR18_14_SIG, ADDR18_15_SIG,
       ADDR18_16_SIG, ADDR18_17_SIG, ADDR18_18_SIG, ADDR18_19_SIG, ADDR18_20_SIG, ADDR18_21_SIG, ADDR18_22_SIG, ADDR18_23_SIG,
       ADDR18_24_SIG, ADDR18_25_SIG, ADDR18_26_SIG, ADDR18_27_SIG, ADDR18_28_SIG, ADDR18_29_SIG, ADDR18_30_SIG, ADDR18_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR19_0_SIG, ADDR19_1_SIG, ADDR19_2_SIG,  ADDR19_3_SIG,  ADDR19_4_SIG,  ADDR19_5_SIG,  ADDR19_6_SIG,  ADDR19_7_SIG,
       ADDR19_8_SIG, ADDR19_9_SIG, ADDR19_10_SIG, ADDR19_11_SIG, ADDR19_12_SIG, ADDR19_13_SIG, ADDR19_14_SIG, ADDR19_15_SIG,
       ADDR19_16_SIG, ADDR19_17_SIG, ADDR19_18_SIG, ADDR19_19_SIG, ADDR19_20_SIG, ADDR19_21_SIG, ADDR19_22_SIG, ADDR19_23_SIG,
       ADDR19_24_SIG, ADDR19_25_SIG, ADDR19_26_SIG, ADDR19_27_SIG, ADDR19_28_SIG, ADDR19_29_SIG, ADDR19_30_SIG, ADDR19_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR20_0_SIG, ADDR20_1_SIG, ADDR20_2_SIG,  ADDR20_3_SIG,  ADDR20_4_SIG,  ADDR20_5_SIG,  ADDR20_6_SIG, ADDR20_7_SIG,
       ADDR20_8_SIG, ADDR20_9_SIG, ADDR20_10_SIG, ADDR20_11_SIG, ADDR20_12_SIG, ADDR20_13_SIG, ADDR20_14_SIG, ADDR20_15_SIG,
       ADDR20_16_SIG, ADDR20_17_SIG, ADDR20_18_SIG, ADDR20_19_SIG, ADDR20_20_SIG, ADDR20_21_SIG, ADDR20_22_SIG, ADDR20_23_SIG,
       ADDR20_24_SIG, ADDR20_25_SIG, ADDR20_26_SIG, ADDR20_27_SIG, ADDR20_28_SIG, ADDR20_29_SIG, ADDR20_30_SIG, ADDR20_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR21_0_SIG, ADDR21_1_SIG, ADDR21_2_SIG,  ADDR21_3_SIG,  ADDR21_4_SIG,  ADDR21_5_SIG,  ADDR21_6_SIG, ADDR21_7_SIG,
       ADDR21_8_SIG, ADDR21_9_SIG, ADDR21_10_SIG, ADDR21_11_SIG, ADDR21_12_SIG, ADDR21_13_SIG, ADDR21_14_SIG, ADDR21_15_SIG,
       ADDR21_16_SIG, ADDR21_17_SIG, ADDR21_18_SIG, ADDR21_19_SIG, ADDR21_20_SIG, ADDR21_21_SIG, ADDR21_22_SIG, ADDR21_23_SIG,
       ADDR21_24_SIG, ADDR21_25_SIG, ADDR21_26_SIG, ADDR21_27_SIG, ADDR21_28_SIG, ADDR21_29_SIG, ADDR21_30_SIG, ADDR21_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR22_0_SIG, ADDR22_1_SIG, ADDR22_2_SIG,  ADDR22_3_SIG,  ADDR22_4_SIG,  ADDR22_5_SIG,  ADDR22_6_SIG,  ADDR22_7_SIG,
       ADDR22_8_SIG, ADDR22_9_SIG, ADDR22_10_SIG, ADDR22_11_SIG, ADDR22_12_SIG, ADDR22_13_SIG, ADDR22_14_SIG, ADDR22_15_SIG,
       ADDR22_16_SIG, ADDR22_17_SIG, ADDR22_18_SIG, ADDR22_19_SIG, ADDR22_20_SIG, ADDR22_21_SIG, ADDR22_22_SIG, ADDR22_23_SIG,
       ADDR22_24_SIG, ADDR22_25_SIG, ADDR22_26_SIG, ADDR22_27_SIG, ADDR22_28_SIG, ADDR22_29_SIG, ADDR22_30_SIG, ADDR22_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR23_0_SIG, ADDR23_1_SIG, ADDR23_2_SIG,  ADDR23_3_SIG, ADDR23_4_SIG,  ADDR23_5_SIG,  ADDR23_6_SIG,  ADDR23_7_SIG,
       ADDR23_8_SIG, ADDR23_9_SIG, ADDR23_10_SIG, ADDR23_11_SIG, ADDR23_12_SIG, ADDR23_13_SIG, ADDR23_14_SIG, ADDR23_15_SIG,
       ADDR23_16_SIG, ADDR23_17_SIG, ADDR23_18_SIG, ADDR23_19_SIG, ADDR23_20_SIG, ADDR23_21_SIG, ADDR23_22_SIG, ADDR23_23_SIG,
       ADDR23_24_SIG, ADDR23_25_SIG, ADDR23_26_SIG, ADDR23_27_SIG, ADDR23_28_SIG, ADDR23_29_SIG, ADDR23_30_SIG, ADDR23_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR24_0_SIG, ADDR24_1_SIG, ADDR24_2_SIG,  ADDR24_3_SIG,  ADDR24_4_SIG,  ADDR24_5_SIG,  ADDR24_6_SIG,  ADDR24_7_SIG,
       ADDR24_8_SIG, ADDR24_9_SIG, ADDR24_10_SIG, ADDR24_11_SIG, ADDR24_12_SIG, ADDR24_13_SIG, ADDR24_14_SIG, ADDR24_15_SIG,
       ADDR24_16_SIG, ADDR24_17_SIG, ADDR24_18_SIG, ADDR24_19_SIG, ADDR24_20_SIG, ADDR24_21_SIG, ADDR24_22_SIG, ADDR24_23_SIG,
       ADDR24_24_SIG, ADDR24_25_SIG, ADDR24_26_SIG, ADDR24_27_SIG, ADDR24_28_SIG, ADDR24_29_SIG, ADDR24_30_SIG, ADDR24_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR25_0_SIG, ADDR25_1_SIG, ADDR25_2_SIG,  ADDR25_3_SIG,  ADDR25_4_SIG,  ADDR25_5_SIG,  ADDR25_6_SIG,  ADDR25_7_SIG,
       ADDR25_8_SIG, ADDR25_9_SIG, ADDR25_10_SIG, ADDR25_11_SIG, ADDR25_12_SIG, ADDR25_13_SIG, ADDR25_14_SIG, ADDR25_15_SIG,
       ADDR25_16_SIG, ADDR25_17_SIG, ADDR25_18_SIG, ADDR25_19_SIG, ADDR25_20_SIG, ADDR25_21_SIG, ADDR25_22_SIG, ADDR25_23_SIG,
       ADDR25_24_SIG, ADDR25_25_SIG, ADDR25_26_SIG, ADDR25_27_SIG, ADDR25_28_SIG, ADDR25_29_SIG, ADDR25_30_SIG, ADDR25_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR26_0_SIG, ADDR26_1_SIG, ADDR26_2_SIG,  ADDR26_3_SIG,  ADDR26_4_SIG,  ADDR26_5_SIG,  ADDR26_6_SIG,  ADDR26_7_SIG,
       ADDR26_8_SIG, ADDR26_9_SIG, ADDR26_10_SIG, ADDR26_11_SIG, ADDR26_12_SIG, ADDR26_13_SIG, ADDR26_14_SIG, ADDR26_15_SIG,
       ADDR26_16_SIG, ADDR26_17_SIG, ADDR26_18_SIG, ADDR26_19_SIG, ADDR26_20_SIG, ADDR26_21_SIG, ADDR26_22_SIG, ADDR26_23_SIG,
       ADDR26_24_SIG, ADDR26_25_SIG, ADDR26_26_SIG, ADDR26_27_SIG, ADDR26_28_SIG, ADDR26_29_SIG, ADDR26_30_SIG, ADDR26_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR27_0_SIG, ADDR27_1_SIG, ADDR27_2_SIG, ADDR27_3_SIG,  ADDR27_4_SIG,  ADDR27_5_SIG,  ADDR27_6_SIG,  ADDR27_7_SIG,
       ADDR27_8_SIG, ADDR27_9_SIG, ADDR27_10_SIG, ADDR27_11_SIG, ADDR27_12_SIG, ADDR27_13_SIG, ADDR27_14_SIG, ADDR27_15_SIG,
       ADDR27_16_SIG, ADDR27_17_SIG, ADDR27_18_SIG, ADDR27_19_SIG, ADDR27_20_SIG, ADDR27_21_SIG, ADDR27_22_SIG, ADDR27_23_SIG,
       ADDR27_24_SIG, ADDR27_25_SIG, ADDR27_26_SIG, ADDR27_27_SIG, ADDR27_28_SIG, ADDR27_29_SIG, ADDR27_30_SIG, ADDR27_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR28_0_SIG, ADDR28_1_SIG, ADDR28_2_SIG,  ADDR28_3_SIG,  ADDR28_4_SIG,  ADDR28_5_SIG,  ADDR28_6_SIG,  ADDR28_7_SIG,
       ADDR28_8_SIG, ADDR28_9_SIG, ADDR28_10_SIG, ADDR28_11_SIG, ADDR28_12_SIG, ADDR28_13_SIG, ADDR28_14_SIG, ADDR28_15_SIG,
       ADDR28_16_SIG, ADDR28_17_SIG, ADDR28_18_SIG, ADDR28_19_SIG, ADDR28_20_SIG, ADDR28_21_SIG, ADDR28_22_SIG, ADDR28_23_SIG,
       ADDR28_24_SIG, ADDR28_25_SIG, ADDR28_26_SIG, ADDR28_27_SIG, ADDR28_28_SIG, ADDR28_29_SIG, ADDR28_30_SIG, ADDR28_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR29_0_SIG, ADDR29_1_SIG, ADDR29_2_SIG,  ADDR29_3_SIG,  ADDR29_4_SIG,  ADDR29_5_SIG,  ADDR29_6_SIG,  ADDR29_7_SIG,
       ADDR29_8_SIG, ADDR29_9_SIG, ADDR29_10_SIG, ADDR29_11_SIG, ADDR29_12_SIG, ADDR29_13_SIG, ADDR29_14_SIG, ADDR29_15_SIG,
       ADDR29_16_SIG, ADDR29_17_SIG, ADDR29_18_SIG, ADDR29_19_SIG, ADDR29_20_SIG, ADDR29_21_SIG, ADDR29_22_SIG, ADDR29_23_SIG,
       ADDR29_24_SIG, ADDR29_25_SIG, ADDR29_26_SIG, ADDR29_27_SIG, ADDR29_28_SIG, ADDR29_29_SIG, ADDR29_30_SIG, ADDR29_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR30_0_SIG, ADDR30_1_SIG, ADDR30_2_SIG,  ADDR30_3_SIG,  ADDR30_4_SIG,  ADDR30_5_SIG,  ADDR30_6_SIG,  ADDR30_7_SIG,
       ADDR30_8_SIG, ADDR30_9_SIG, ADDR30_10_SIG, ADDR30_11_SIG, ADDR30_12_SIG, ADDR30_13_SIG, ADDR30_14_SIG, ADDR30_15_SIG,
       ADDR30_16_SIG, ADDR30_17_SIG, ADDR30_18_SIG, ADDR30_19_SIG, ADDR30_20_SIG, ADDR30_21_SIG, ADDR30_22_SIG, ADDR30_23_SIG,
       ADDR30_24_SIG, ADDR30_25_SIG, ADDR30_26_SIG, ADDR30_27_SIG, ADDR30_28_SIG, ADDR30_29_SIG, ADDR30_30_SIG, ADDR30_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal ADDR31_0_SIG, ADDR31_1_SIG, ADDR31_2_SIG,  ADDR31_3_SIG,  ADDR31_4_SIG,  ADDR31_5_SIG,  ADDR31_6_SIG,  ADDR31_7_SIG,
       ADDR31_8_SIG, ADDR31_9_SIG, ADDR31_10_SIG, ADDR31_11_SIG, ADDR31_12_SIG, ADDR31_13_SIG, ADDR31_14_SIG, ADDR31_15_SIG,
       ADDR31_16_SIG, ADDR31_17_SIG, ADDR31_18_SIG, ADDR31_19_SIG, ADDR31_20_SIG, ADDR31_21_SIG, ADDR31_22_SIG, ADDR31_23_SIG,
       ADDR31_24_SIG, ADDR31_25_SIG, ADDR31_26_SIG, ADDR31_27_SIG, ADDR31_28_SIG, ADDR31_29_SIG, ADDR31_30_SIG, ADDR31_31_SIG : std_logic_vector(POWER-1 downto 0):= (others => '0');
signal BIAS0_ROM_ADDR  : std_logic_vector(4 downto 0) := "00000";
signal BIAS1_ROM_ADDR  : std_logic_vector(4 downto 0) := "00001";
signal BIAS2_ROM_ADDR  : std_logic_vector(4 downto 0) := "00010";
signal BIAS3_ROM_ADDR  : std_logic_vector(4 downto 0) := "00011";
signal BIAS4_ROM_ADDR  : std_logic_vector(4 downto 0) := "00100";
signal BIAS5_ROM_ADDR  : std_logic_vector(4 downto 0) := "00101";
signal BIAS6_ROM_ADDR  : std_logic_vector(4 downto 0) := "00110";
signal BIAS7_ROM_ADDR  : std_logic_vector(4 downto 0) := "00111";
signal BIAS8_ROM_ADDR  : std_logic_vector(4 downto 0) := "01000";
signal BIAS9_ROM_ADDR  : std_logic_vector(4 downto 0) := "01001";
signal BIAS10_ROM_ADDR : std_logic_vector(4 downto 0) := "01010";
signal BIAS11_ROM_ADDR : std_logic_vector(4 downto 0) := "01011";
signal BIAS12_ROM_ADDR : std_logic_vector(4 downto 0) := "01100";
signal BIAS13_ROM_ADDR : std_logic_vector(4 downto 0) := "01101";
signal BIAS14_ROM_ADDR : std_logic_vector(4 downto 0) := "01110";
signal BIAS15_ROM_ADDR : std_logic_vector(4 downto 0) := "01111";
signal BIAS16_ROM_ADDR : std_logic_vector(4 downto 0) := "10000";
signal BIAS17_ROM_ADDR : std_logic_vector(4 downto 0) := "10001";
signal BIAS18_ROM_ADDR : std_logic_vector(4 downto 0) := "10010";
signal BIAS19_ROM_ADDR : std_logic_vector(4 downto 0) := "10011";
signal BIAS20_ROM_ADDR : std_logic_vector(4 downto 0) := "10100";
signal BIAS21_ROM_ADDR : std_logic_vector(4 downto 0) := "10101";
signal BIAS22_ROM_ADDR : std_logic_vector(4 downto 0) := "10110";
signal BIAS23_ROM_ADDR : std_logic_vector(4 downto 0) := "10111";
signal BIAS24_ROM_ADDR : std_logic_vector(4 downto 0) := "11000";
signal BIAS25_ROM_ADDR : std_logic_vector(4 downto 0) := "11001";
signal BIAS26_ROM_ADDR : std_logic_vector(4 downto 0) := "11010";
signal BIAS27_ROM_ADDR : std_logic_vector(4 downto 0) := "11011";
signal BIAS28_ROM_ADDR : std_logic_vector(4 downto 0) := "11100";
signal BIAS29_ROM_ADDR : std_logic_vector(4 downto 0) := "11101"; 
signal BIAS0_SIG, BIAS1_SIG, BIAS2_SIG, BIAS3_SIG, BIAS4_SIG,
       BIAS5_SIG, BIAS6_SIG, BIAS7_SIG, BIAS8_SIG, BIAS9_SIG,
       BIAS10_SIG, BIAS11_SIG, BIAS12_SIG, BIAS13_SIG, BIAS14_SIG,
       BIAS15_SIG, BIAS16_SIG, BIAS17_SIG, BIAS18_SIG, BIAS19_SIG,
       BIAS20_SIG, BIAS21_SIG, BIAS22_SIG, BIAS23_SIG, BIAS24_SIG,
       BIAS25_SIG, BIAS26_SIG, BIAS27_SIG, BIAS28_SIG, BIAS29_SIG : std_logic_vector(WIDTH+WIDTH-1 downto 0) := (others => '0');
signal VM0_OUT_SIG, VM1_OUT_SIG, VM2_OUT_SIG, VM3_OUT_SIG, VM4_OUT_SIG,
       VM5_OUT_SIG, VM6_OUT_SIG, VM7_OUT_SIG, VM8_OUT_SIG, VM9_OUT_SIG,
       VM10_OUT_SIG, VM11_OUT_SIG, VM12_OUT_SIG, VM13_OUT_SIG, VM14_OUT_SIG,
       VM15_OUT_SIG, VM16_OUT_SIG, VM17_OUT_SIG, VM18_OUT_SIG, VM19_OUT_SIG,
       VM20_OUT_SIG, VM21_OUT_SIG, VM22_OUT_SIG, VM23_OUT_SIG, VM24_OUT_SIG,
       VM25_OUT_SIG, VM26_OUT_SIG, VM27_OUT_SIG, VM28_OUT_SIG, VM29_OUT_SIG  :  std_logic_vector(WIDTH+WIDTH-1 downto 0) := (others => '0');
signal ADDER0_OUT_SIG, ADDER1_OUT_SIG, ADDER2_OUT_SIG, ADDER3_OUT_SIG, ADDER4_OUT_SIG,
       ADDER5_OUT_SIG, ADDER6_OUT_SIG, ADDER7_OUT_SIG, ADDER8_OUT_SIG, ADDER9_OUT_SIG,
       ADDER10_OUT_SIG, ADDER11_OUT_SIG, ADDER12_OUT_SIG, ADDER13_OUT_SIG, ADDER14_OUT_SIG,
       ADDER15_OUT_SIG, ADDER16_OUT_SIG, ADDER17_OUT_SIG, ADDER18_OUT_SIG, ADDER19_OUT_SIG,
       ADDER20_OUT_SIG, ADDER21_OUT_SIG, ADDER22_OUT_SIG, ADDER23_OUT_SIG, ADDER24_OUT_SIG,
       ADDER25_OUT_SIG, ADDER26_OUT_SIG, ADDER27_OUT_SIG, ADDER28_OUT_SIG, ADDER29_OUT_SIG : std_logic_vector(WIDTH+WIDTH-1 downto 0) := (others => '0');
signal SET_VM_SIG, SET_CNT_SIG: std_logic := '0';

begin

SET_CNT_SIG <= SET_CNT; 

DIN0_SIG  <= DIN0;
DIN1_SIG  <= DIN1;
DIN2_SIG  <= DIN2;
DIN3_SIG  <= DIN3;
DIN4_SIG  <= DIN4;
DIN5_SIG  <= DIN5;
DIN6_SIG  <= DIN6;
DIN7_SIG  <= DIN7;
DIN8_SIG  <= DIN8;
DIN9_SIG  <= DIN9;
DIN10_SIG  <= DIN10;
DIN11_SIG  <= DIN11;
DIN12_SIG  <= DIN12;
DIN13_SIG  <= DIN13;
DIN14_SIG  <= DIN14;
DIN15_SIG  <= DIN15;
DIN16_SIG  <= DIN16;
DIN17_SIG  <= DIN17;
DIN18_SIG  <= DIN18;
DIN19_SIG  <= DIN19;
DIN20_SIG  <= DIN20;
DIN21_SIG  <= DIN21;
DIN22_SIG  <= DIN22;
DIN23_SIG  <= DIN23;
DIN24_SIG  <= DIN24;
DIN25_SIG  <= DIN25;
DIN26_SIG  <= DIN26;
DIN27_SIG  <= DIN27;
DIN28_SIG  <= DIN28;
DIN29_SIG  <= DIN29;
DIN30_SIG  <= DIN30;
DIN31_SIG  <= DIN31;

VM0_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM0_DATA0_SIG,
    ROM1_DATA   => ROM0_DATA1_SIG,
    ROM2_DATA   => ROM0_DATA2_SIG,
    ROM3_DATA   => ROM0_DATA3_SIG,
    ROM4_DATA   => ROM0_DATA4_SIG,
    ROM5_DATA   => ROM0_DATA5_SIG,
    ROM6_DATA   => ROM0_DATA6_SIG,
    ROM7_DATA   => ROM0_DATA7_SIG,
    ROM8_DATA   => ROM0_DATA8_SIG,
    ROM9_DATA   => ROM0_DATA9_SIG,
    ROM10_DATA  => ROM0_DATA10_SIG,
    ROM11_DATA  => ROM0_DATA11_SIG,
    ROM12_DATA  => ROM0_DATA12_SIG,
    ROM13_DATA  => ROM0_DATA13_SIG,
    ROM14_DATA  => ROM0_DATA14_SIG,
    ROM15_DATA  => ROM0_DATA15_SIG,
    ROM16_DATA  => ROM0_DATA16_SIG,
    ROM17_DATA  => ROM0_DATA17_SIG,
    ROM18_DATA  => ROM0_DATA18_SIG,
    ROM19_DATA  => ROM0_DATA19_SIG,
    ROM20_DATA  => ROM0_DATA20_SIG,
    ROM21_DATA  => ROM0_DATA21_SIG,
    ROM22_DATA  => ROM0_DATA22_SIG,
    ROM23_DATA  => ROM0_DATA23_SIG,
    ROM24_DATA  => ROM0_DATA24_SIG,
    ROM25_DATA  => ROM0_DATA25_SIG,
    ROM26_DATA  => ROM0_DATA26_SIG,
    ROM27_DATA  => ROM0_DATA27_SIG,
    ROM28_DATA  => ROM0_DATA28_SIG,
    ROM29_DATA  => ROM0_DATA29_SIG,
    ROM30_DATA  => ROM0_DATA30_SIG,
    ROM31_DATA  => ROM0_DATA31_SIG,
    ADDR0       => ADDR0_0_SIG,
    ADDR1       => ADDR0_1_SIG,
    ADDR2       => ADDR0_2_SIG,
    ADDR3       => ADDR0_3_SIG,
    ADDR4       => ADDR0_4_SIG,
    ADDR5       => ADDR0_5_SIG,
    ADDR6       => ADDR0_6_SIG,
    ADDR7       => ADDR0_7_SIG,
    ADDR8       => ADDR0_8_SIG,
    ADDR9       => ADDR0_9_SIG,
    ADDR10      => ADDR0_10_SIG,
    ADDR11      => ADDR0_11_SIG,
    ADDR12      => ADDR0_12_SIG,
    ADDR13      => ADDR0_13_SIG,
    ADDR14      => ADDR0_14_SIG,
    ADDR15      => ADDR0_15_SIG,
    ADDR16      => ADDR0_16_SIG,
    ADDR17      => ADDR0_17_SIG,
    ADDR18      => ADDR0_18_SIG,
    ADDR19      => ADDR0_19_SIG,
    ADDR20      => ADDR0_20_SIG,
    ADDR21      => ADDR0_21_SIG,
    ADDR22      => ADDR0_22_SIG,
    ADDR23      => ADDR0_23_SIG,
    ADDR24      => ADDR0_24_SIG,
    ADDR25      => ADDR0_25_SIG,
    ADDR26      => ADDR0_26_SIG,
    ADDR27      => ADDR0_27_SIG,
    ADDR28      => ADDR0_28_SIG,
    ADDR29      => ADDR0_29_SIG,
    ADDR30      => ADDR0_30_SIG,
    ADDR31      => ADDR0_31_SIG,
    DOUT        => VM0_OUT_SIG
);

VM1_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM1_DATA0_SIG,
    ROM1_DATA   => ROM1_DATA1_SIG,
    ROM2_DATA   => ROM1_DATA2_SIG,
    ROM3_DATA   => ROM1_DATA3_SIG,
    ROM4_DATA   => ROM1_DATA4_SIG,
    ROM5_DATA   => ROM1_DATA5_SIG,
    ROM6_DATA   => ROM1_DATA6_SIG,
    ROM7_DATA   => ROM1_DATA7_SIG,
    ROM8_DATA   => ROM1_DATA8_SIG,
    ROM9_DATA   => ROM1_DATA9_SIG,
    ROM10_DATA  => ROM1_DATA10_SIG,
    ROM11_DATA  => ROM1_DATA11_SIG,
    ROM12_DATA  => ROM1_DATA12_SIG,
    ROM13_DATA  => ROM1_DATA13_SIG,
    ROM14_DATA  => ROM1_DATA14_SIG,
    ROM15_DATA  => ROM1_DATA15_SIG,
    ROM16_DATA  => ROM1_DATA16_SIG,
    ROM17_DATA  => ROM1_DATA17_SIG,
    ROM18_DATA  => ROM1_DATA18_SIG,
    ROM19_DATA  => ROM1_DATA19_SIG,
    ROM20_DATA  => ROM1_DATA20_SIG,
    ROM21_DATA  => ROM1_DATA21_SIG,
    ROM22_DATA  => ROM1_DATA22_SIG,
    ROM23_DATA  => ROM1_DATA23_SIG,
    ROM24_DATA  => ROM1_DATA24_SIG,
    ROM25_DATA  => ROM1_DATA25_SIG,
    ROM26_DATA  => ROM1_DATA26_SIG,
    ROM27_DATA  => ROM1_DATA27_SIG,
    ROM28_DATA  => ROM1_DATA28_SIG,
    ROM29_DATA  => ROM1_DATA29_SIG,
    ROM30_DATA  => ROM1_DATA30_SIG,
    ROM31_DATA  => ROM1_DATA31_SIG,
    ADDR0       => ADDR1_0_SIG,
    ADDR1       => ADDR1_1_SIG,
    ADDR2       => ADDR1_2_SIG,
    ADDR3       => ADDR1_3_SIG,
    ADDR4       => ADDR1_4_SIG,
    ADDR5       => ADDR1_5_SIG,
    ADDR6       => ADDR1_6_SIG,
    ADDR7       => ADDR1_7_SIG,
    ADDR8       => ADDR1_8_SIG,
    ADDR9       => ADDR1_9_SIG,
    ADDR10      => ADDR1_10_SIG,
    ADDR11      => ADDR1_11_SIG,
    ADDR12      => ADDR1_12_SIG,
    ADDR13      => ADDR1_13_SIG,
    ADDR14      => ADDR1_14_SIG,
    ADDR15      => ADDR1_15_SIG,
    ADDR16      => ADDR1_16_SIG,
    ADDR17      => ADDR1_17_SIG,
    ADDR18      => ADDR1_18_SIG,
    ADDR19      => ADDR1_19_SIG,
    ADDR20      => ADDR1_20_SIG,
    ADDR21      => ADDR1_21_SIG,
    ADDR22      => ADDR1_22_SIG,
    ADDR23      => ADDR1_23_SIG,
    ADDR24      => ADDR1_24_SIG,
    ADDR25      => ADDR1_25_SIG,
    ADDR26      => ADDR1_26_SIG,
    ADDR27      => ADDR1_27_SIG,
    ADDR28      => ADDR1_28_SIG,
    ADDR29      => ADDR1_29_SIG,
    ADDR30      => ADDR1_30_SIG,
    ADDR31      => ADDR1_31_SIG,
    DOUT        => VM1_OUT_SIG
);

VM2_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM2_DATA0_SIG,
    ROM1_DATA   => ROM2_DATA1_SIG,
    ROM2_DATA   => ROM2_DATA2_SIG,
    ROM3_DATA   => ROM2_DATA3_SIG,
    ROM4_DATA   => ROM2_DATA4_SIG,
    ROM5_DATA   => ROM2_DATA5_SIG,
    ROM6_DATA   => ROM2_DATA6_SIG,
    ROM7_DATA   => ROM2_DATA7_SIG,
    ROM8_DATA   => ROM2_DATA8_SIG,
    ROM9_DATA   => ROM2_DATA9_SIG,
    ROM10_DATA  => ROM2_DATA10_SIG,
    ROM11_DATA  => ROM2_DATA11_SIG,
    ROM12_DATA  => ROM2_DATA12_SIG,
    ROM13_DATA  => ROM2_DATA13_SIG,
    ROM14_DATA  => ROM2_DATA14_SIG,
    ROM15_DATA  => ROM2_DATA15_SIG,
    ROM16_DATA  => ROM2_DATA16_SIG,
    ROM17_DATA  => ROM2_DATA17_SIG,
    ROM18_DATA  => ROM2_DATA18_SIG,
    ROM19_DATA  => ROM2_DATA19_SIG,
    ROM20_DATA  => ROM2_DATA20_SIG,
    ROM21_DATA  => ROM2_DATA21_SIG,
    ROM22_DATA  => ROM2_DATA22_SIG,
    ROM23_DATA  => ROM2_DATA23_SIG,
    ROM24_DATA  => ROM2_DATA24_SIG,
    ROM25_DATA  => ROM2_DATA25_SIG,
    ROM26_DATA  => ROM2_DATA26_SIG,
    ROM27_DATA  => ROM2_DATA27_SIG,
    ROM28_DATA  => ROM2_DATA28_SIG,
    ROM29_DATA  => ROM2_DATA29_SIG,
    ROM30_DATA  => ROM2_DATA30_SIG,
    ROM31_DATA  => ROM2_DATA31_SIG,
    ADDR0       => ADDR2_0_SIG,
    ADDR1       => ADDR2_1_SIG,
    ADDR2       => ADDR2_2_SIG,
    ADDR3       => ADDR2_3_SIG,
    ADDR4       => ADDR2_4_SIG,
    ADDR5       => ADDR2_5_SIG,
    ADDR6       => ADDR2_6_SIG,
    ADDR7       => ADDR2_7_SIG,
    ADDR8       => ADDR2_8_SIG,
    ADDR9       => ADDR2_9_SIG,
    ADDR10      => ADDR2_10_SIG,
    ADDR11      => ADDR2_11_SIG,
    ADDR12      => ADDR2_12_SIG,
    ADDR13      => ADDR2_13_SIG,
    ADDR14      => ADDR2_14_SIG,
    ADDR15      => ADDR2_15_SIG,
    ADDR16      => ADDR2_16_SIG,
    ADDR17      => ADDR2_17_SIG,
    ADDR18      => ADDR2_18_SIG,
    ADDR19      => ADDR2_19_SIG,
    ADDR20      => ADDR2_20_SIG,
    ADDR21      => ADDR2_21_SIG,
    ADDR22      => ADDR2_22_SIG,
    ADDR23      => ADDR2_23_SIG,
    ADDR24      => ADDR2_24_SIG,
    ADDR25      => ADDR2_25_SIG,
    ADDR26      => ADDR2_26_SIG,
    ADDR27      => ADDR2_27_SIG,
    ADDR28      => ADDR2_28_SIG,
    ADDR29      => ADDR2_29_SIG,
    ADDR30      => ADDR2_30_SIG,
    ADDR31      => ADDR2_31_SIG,
    DOUT        => VM2_OUT_SIG
);

VM3_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM3_DATA0_SIG,
    ROM1_DATA   => ROM3_DATA1_SIG,
    ROM2_DATA   => ROM3_DATA2_SIG,
    ROM3_DATA   => ROM3_DATA3_SIG,
    ROM4_DATA   => ROM3_DATA4_SIG,
    ROM5_DATA   => ROM3_DATA5_SIG,
    ROM6_DATA   => ROM3_DATA6_SIG,
    ROM7_DATA   => ROM3_DATA7_SIG,
    ROM8_DATA   => ROM3_DATA8_SIG,
    ROM9_DATA   => ROM3_DATA9_SIG,
    ROM10_DATA  => ROM3_DATA10_SIG,
    ROM11_DATA  => ROM3_DATA11_SIG,
    ROM12_DATA  => ROM3_DATA12_SIG,
    ROM13_DATA  => ROM3_DATA13_SIG,
    ROM14_DATA  => ROM3_DATA14_SIG,
    ROM15_DATA  => ROM3_DATA15_SIG,
    ROM16_DATA  => ROM3_DATA16_SIG,
    ROM17_DATA  => ROM3_DATA17_SIG,
    ROM18_DATA  => ROM3_DATA18_SIG,
    ROM19_DATA  => ROM3_DATA19_SIG,
    ROM20_DATA  => ROM3_DATA20_SIG,
    ROM21_DATA  => ROM3_DATA21_SIG,
    ROM22_DATA  => ROM3_DATA22_SIG,
    ROM23_DATA  => ROM3_DATA23_SIG,
    ROM24_DATA  => ROM3_DATA24_SIG,
    ROM25_DATA  => ROM3_DATA25_SIG,
    ROM26_DATA  => ROM3_DATA26_SIG,
    ROM27_DATA  => ROM3_DATA27_SIG,
    ROM28_DATA  => ROM3_DATA28_SIG,
    ROM29_DATA  => ROM3_DATA29_SIG,
    ROM30_DATA  => ROM3_DATA30_SIG,
    ROM31_DATA  => ROM3_DATA31_SIG,
    ADDR0       => ADDR3_0_SIG,
    ADDR1       => ADDR3_1_SIG,
    ADDR2       => ADDR3_2_SIG,
    ADDR3       => ADDR3_3_SIG,
    ADDR4       => ADDR3_4_SIG,
    ADDR5       => ADDR3_5_SIG,
    ADDR6       => ADDR3_6_SIG,
    ADDR7       => ADDR3_7_SIG,
    ADDR8       => ADDR3_8_SIG,
    ADDR9       => ADDR3_9_SIG,
    ADDR10      => ADDR3_10_SIG,
    ADDR11      => ADDR3_11_SIG,
    ADDR12      => ADDR3_12_SIG,
    ADDR13      => ADDR3_13_SIG,
    ADDR14      => ADDR3_14_SIG,
    ADDR15      => ADDR3_15_SIG,
    ADDR16      => ADDR3_16_SIG,
    ADDR17      => ADDR3_17_SIG,
    ADDR18      => ADDR3_18_SIG,
    ADDR19      => ADDR3_19_SIG,
    ADDR20      => ADDR3_20_SIG,
    ADDR21      => ADDR3_21_SIG,
    ADDR22      => ADDR3_22_SIG,
    ADDR23      => ADDR3_23_SIG,
    ADDR24      => ADDR3_24_SIG,
    ADDR25      => ADDR3_25_SIG,
    ADDR26      => ADDR3_26_SIG,
    ADDR27      => ADDR3_27_SIG,
    ADDR28      => ADDR3_28_SIG,
    ADDR29      => ADDR3_29_SIG,
    ADDR30      => ADDR3_30_SIG,
    ADDR31      => ADDR3_31_SIG,
    DOUT        => VM3_OUT_SIG
);

VM4_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM4_DATA0_SIG,
    ROM1_DATA   => ROM4_DATA1_SIG,
    ROM2_DATA   => ROM4_DATA2_SIG,
    ROM3_DATA   => ROM4_DATA3_SIG,
    ROM4_DATA   => ROM4_DATA4_SIG,
    ROM5_DATA   => ROM4_DATA5_SIG,
    ROM6_DATA   => ROM4_DATA6_SIG,
    ROM7_DATA   => ROM4_DATA7_SIG,
    ROM8_DATA   => ROM4_DATA8_SIG,
    ROM9_DATA   => ROM4_DATA9_SIG,
    ROM10_DATA  => ROM4_DATA10_SIG,
    ROM11_DATA  => ROM4_DATA11_SIG,
    ROM12_DATA  => ROM4_DATA12_SIG,
    ROM13_DATA  => ROM4_DATA13_SIG,
    ROM14_DATA  => ROM4_DATA14_SIG,
    ROM15_DATA  => ROM4_DATA15_SIG,
    ROM16_DATA  => ROM4_DATA16_SIG,
    ROM17_DATA  => ROM4_DATA17_SIG,
    ROM18_DATA  => ROM4_DATA18_SIG,
    ROM19_DATA  => ROM4_DATA19_SIG,
    ROM20_DATA  => ROM4_DATA20_SIG,
    ROM21_DATA  => ROM4_DATA21_SIG,
    ROM22_DATA  => ROM4_DATA22_SIG,
    ROM23_DATA  => ROM4_DATA23_SIG,
    ROM24_DATA  => ROM4_DATA24_SIG,
    ROM25_DATA  => ROM4_DATA25_SIG,
    ROM26_DATA  => ROM4_DATA26_SIG,
    ROM27_DATA  => ROM4_DATA27_SIG,
    ROM28_DATA  => ROM4_DATA28_SIG,
    ROM29_DATA  => ROM4_DATA29_SIG,
    ROM30_DATA  => ROM4_DATA30_SIG,
    ROM31_DATA  => ROM4_DATA31_SIG,
    ADDR0       => ADDR4_0_SIG,
    ADDR1       => ADDR4_1_SIG,
    ADDR2       => ADDR4_2_SIG,
    ADDR3       => ADDR4_3_SIG,
    ADDR4       => ADDR4_4_SIG,
    ADDR5       => ADDR4_5_SIG,
    ADDR6       => ADDR4_6_SIG,
    ADDR7       => ADDR4_7_SIG,
    ADDR8       => ADDR4_8_SIG,
    ADDR9       => ADDR4_9_SIG,
    ADDR10      => ADDR4_10_SIG,
    ADDR11      => ADDR4_11_SIG,
    ADDR12      => ADDR4_12_SIG,
    ADDR13      => ADDR4_13_SIG,
    ADDR14      => ADDR4_14_SIG,
    ADDR15      => ADDR4_15_SIG,
    ADDR16      => ADDR4_16_SIG,
    ADDR17      => ADDR4_17_SIG,
    ADDR18      => ADDR4_18_SIG,
    ADDR19      => ADDR4_19_SIG,
    ADDR20      => ADDR4_20_SIG,
    ADDR21      => ADDR4_21_SIG,
    ADDR22      => ADDR4_22_SIG,
    ADDR23      => ADDR4_23_SIG,
    ADDR24      => ADDR4_24_SIG,
    ADDR25      => ADDR4_25_SIG,
    ADDR26      => ADDR4_26_SIG,
    ADDR27      => ADDR4_27_SIG,
    ADDR28      => ADDR4_28_SIG,
    ADDR29      => ADDR4_29_SIG,
    ADDR30      => ADDR4_30_SIG,
    ADDR31      => ADDR4_31_SIG,
    DOUT        => VM4_OUT_SIG
);

VM5_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM5_DATA0_SIG,
    ROM1_DATA   => ROM5_DATA1_SIG,
    ROM2_DATA   => ROM5_DATA2_SIG,
    ROM3_DATA   => ROM5_DATA3_SIG,
    ROM4_DATA   => ROM5_DATA4_SIG,
    ROM5_DATA   => ROM5_DATA5_SIG,
    ROM6_DATA   => ROM5_DATA6_SIG,
    ROM7_DATA   => ROM5_DATA7_SIG,
    ROM8_DATA   => ROM5_DATA8_SIG,
    ROM9_DATA   => ROM5_DATA9_SIG,
    ROM10_DATA  => ROM5_DATA10_SIG,
    ROM11_DATA  => ROM5_DATA11_SIG,
    ROM12_DATA  => ROM5_DATA12_SIG,
    ROM13_DATA  => ROM5_DATA13_SIG,
    ROM14_DATA  => ROM5_DATA14_SIG,
    ROM15_DATA  => ROM5_DATA15_SIG,
    ROM16_DATA  => ROM5_DATA16_SIG,
    ROM17_DATA  => ROM5_DATA17_SIG,
    ROM18_DATA  => ROM5_DATA18_SIG,
    ROM19_DATA  => ROM5_DATA19_SIG,
    ROM20_DATA  => ROM5_DATA20_SIG,
    ROM21_DATA  => ROM5_DATA21_SIG,
    ROM22_DATA  => ROM5_DATA22_SIG,
    ROM23_DATA  => ROM5_DATA23_SIG,
    ROM24_DATA  => ROM5_DATA24_SIG,
    ROM25_DATA  => ROM5_DATA25_SIG,
    ROM26_DATA  => ROM5_DATA26_SIG,
    ROM27_DATA  => ROM5_DATA27_SIG,
    ROM28_DATA  => ROM5_DATA28_SIG,
    ROM29_DATA  => ROM5_DATA29_SIG,
    ROM30_DATA  => ROM5_DATA30_SIG,
    ROM31_DATA  => ROM5_DATA31_SIG,
    ADDR0       => ADDR5_0_SIG,
    ADDR1       => ADDR5_1_SIG,
    ADDR2       => ADDR5_2_SIG,
    ADDR3       => ADDR5_3_SIG,
    ADDR4       => ADDR5_4_SIG,
    ADDR5       => ADDR5_5_SIG,
    ADDR6       => ADDR5_6_SIG,
    ADDR7       => ADDR5_7_SIG,
    ADDR8       => ADDR5_8_SIG,
    ADDR9       => ADDR5_9_SIG,
    ADDR10      => ADDR5_10_SIG,
    ADDR11      => ADDR5_11_SIG,
    ADDR12      => ADDR5_12_SIG,
    ADDR13      => ADDR5_13_SIG,
    ADDR14      => ADDR5_14_SIG,
    ADDR15      => ADDR5_15_SIG,
    ADDR16      => ADDR5_16_SIG,
    ADDR17      => ADDR5_17_SIG,
    ADDR18      => ADDR5_18_SIG,
    ADDR19      => ADDR5_19_SIG,
    ADDR20      => ADDR5_20_SIG,
    ADDR21      => ADDR5_21_SIG,
    ADDR22      => ADDR5_22_SIG,
    ADDR23      => ADDR5_23_SIG,
    ADDR24      => ADDR5_24_SIG,
    ADDR25      => ADDR5_25_SIG,
    ADDR26      => ADDR5_26_SIG,
    ADDR27      => ADDR5_27_SIG,
    ADDR28      => ADDR5_28_SIG,
    ADDR29      => ADDR5_29_SIG,
    ADDR30      => ADDR5_30_SIG,
    ADDR31      => ADDR5_31_SIG,
    DOUT        => VM5_OUT_SIG
);

VM6_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM6_DATA0_SIG,
    ROM1_DATA   => ROM6_DATA1_SIG,
    ROM2_DATA   => ROM6_DATA2_SIG,
    ROM3_DATA   => ROM6_DATA3_SIG,
    ROM4_DATA   => ROM6_DATA4_SIG,
    ROM5_DATA   => ROM6_DATA5_SIG,
    ROM6_DATA   => ROM6_DATA6_SIG,
    ROM7_DATA   => ROM6_DATA7_SIG,
    ROM8_DATA   => ROM6_DATA8_SIG,
    ROM9_DATA   => ROM6_DATA9_SIG,
    ROM10_DATA  => ROM6_DATA10_SIG,
    ROM11_DATA  => ROM6_DATA11_SIG,
    ROM12_DATA  => ROM6_DATA12_SIG,
    ROM13_DATA  => ROM6_DATA13_SIG,
    ROM14_DATA  => ROM6_DATA14_SIG,
    ROM15_DATA  => ROM6_DATA15_SIG,
    ROM16_DATA  => ROM6_DATA16_SIG,
    ROM17_DATA  => ROM6_DATA17_SIG,
    ROM18_DATA  => ROM6_DATA18_SIG,
    ROM19_DATA  => ROM6_DATA19_SIG,
    ROM20_DATA  => ROM6_DATA20_SIG,
    ROM21_DATA  => ROM6_DATA21_SIG,
    ROM22_DATA  => ROM6_DATA22_SIG,
    ROM23_DATA  => ROM6_DATA23_SIG,
    ROM24_DATA  => ROM6_DATA24_SIG,
    ROM25_DATA  => ROM6_DATA25_SIG,
    ROM26_DATA  => ROM6_DATA26_SIG,
    ROM27_DATA  => ROM6_DATA27_SIG,
    ROM28_DATA  => ROM6_DATA28_SIG,
    ROM29_DATA  => ROM6_DATA29_SIG,
    ROM30_DATA  => ROM6_DATA30_SIG,
    ROM31_DATA  => ROM6_DATA31_SIG,
    ADDR0       => ADDR6_0_SIG,
    ADDR1       => ADDR6_1_SIG,
    ADDR2       => ADDR6_2_SIG,
    ADDR3       => ADDR6_3_SIG,
    ADDR4       => ADDR6_4_SIG,
    ADDR5       => ADDR6_5_SIG,
    ADDR6       => ADDR6_6_SIG,
    ADDR7       => ADDR6_7_SIG,
    ADDR8       => ADDR6_8_SIG,
    ADDR9       => ADDR6_9_SIG,
    ADDR10      => ADDR6_10_SIG,
    ADDR11      => ADDR6_11_SIG,
    ADDR12      => ADDR6_12_SIG,
    ADDR13      => ADDR6_13_SIG,
    ADDR14      => ADDR6_14_SIG,
    ADDR15      => ADDR6_15_SIG,
    ADDR16      => ADDR6_16_SIG,
    ADDR17      => ADDR6_17_SIG,
    ADDR18      => ADDR6_18_SIG,
    ADDR19      => ADDR6_19_SIG,
    ADDR20      => ADDR6_20_SIG,
    ADDR21      => ADDR6_21_SIG,
    ADDR22      => ADDR6_22_SIG,
    ADDR23      => ADDR6_23_SIG,
    ADDR24      => ADDR6_24_SIG,
    ADDR25      => ADDR6_25_SIG,
    ADDR26      => ADDR6_26_SIG,
    ADDR27      => ADDR6_27_SIG,
    ADDR28      => ADDR6_28_SIG,
    ADDR29      => ADDR6_29_SIG,
    ADDR30      => ADDR6_30_SIG,
    ADDR31      => ADDR6_31_SIG,
    DOUT        => VM6_OUT_SIG
);

VM7_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM7_DATA0_SIG,
    ROM1_DATA   => ROM7_DATA1_SIG,
    ROM2_DATA   => ROM7_DATA2_SIG,
    ROM3_DATA   => ROM7_DATA3_SIG,
    ROM4_DATA   => ROM7_DATA4_SIG,
    ROM5_DATA   => ROM7_DATA5_SIG,
    ROM6_DATA   => ROM7_DATA6_SIG,
    ROM7_DATA   => ROM7_DATA7_SIG,
    ROM8_DATA   => ROM7_DATA8_SIG,
    ROM9_DATA   => ROM7_DATA9_SIG,
    ROM10_DATA  => ROM7_DATA10_SIG,
    ROM11_DATA  => ROM7_DATA11_SIG,
    ROM12_DATA  => ROM7_DATA12_SIG,
    ROM13_DATA  => ROM7_DATA13_SIG,
    ROM14_DATA  => ROM7_DATA14_SIG,
    ROM15_DATA  => ROM7_DATA15_SIG,
    ROM16_DATA  => ROM7_DATA16_SIG,
    ROM17_DATA  => ROM7_DATA17_SIG,
    ROM18_DATA  => ROM7_DATA18_SIG,
    ROM19_DATA  => ROM7_DATA19_SIG,
    ROM20_DATA  => ROM7_DATA20_SIG,
    ROM21_DATA  => ROM7_DATA21_SIG,
    ROM22_DATA  => ROM7_DATA22_SIG,
    ROM23_DATA  => ROM7_DATA23_SIG,
    ROM24_DATA  => ROM7_DATA24_SIG,
    ROM25_DATA  => ROM7_DATA25_SIG,
    ROM26_DATA  => ROM7_DATA26_SIG,
    ROM27_DATA  => ROM7_DATA27_SIG,
    ROM28_DATA  => ROM7_DATA28_SIG,
    ROM29_DATA  => ROM7_DATA29_SIG,
    ROM30_DATA  => ROM7_DATA30_SIG,
    ROM31_DATA  => ROM7_DATA31_SIG,
    ADDR0       => ADDR7_0_SIG,
    ADDR1       => ADDR7_1_SIG,
    ADDR2       => ADDR7_2_SIG,
    ADDR3       => ADDR7_3_SIG,
    ADDR4       => ADDR7_4_SIG,
    ADDR5       => ADDR7_5_SIG,
    ADDR6       => ADDR7_6_SIG,
    ADDR7       => ADDR7_7_SIG,
    ADDR8       => ADDR7_8_SIG,
    ADDR9       => ADDR7_9_SIG,
    ADDR10      => ADDR7_10_SIG,
    ADDR11      => ADDR7_11_SIG,
    ADDR12      => ADDR7_12_SIG,
    ADDR13      => ADDR7_13_SIG,
    ADDR14      => ADDR7_14_SIG,
    ADDR15      => ADDR7_15_SIG,
    ADDR16      => ADDR7_16_SIG,
    ADDR17      => ADDR7_17_SIG,
    ADDR18      => ADDR7_18_SIG,
    ADDR19      => ADDR7_19_SIG,
    ADDR20      => ADDR7_20_SIG,
    ADDR21      => ADDR7_21_SIG,
    ADDR22      => ADDR7_22_SIG,
    ADDR23      => ADDR7_23_SIG,
    ADDR24      => ADDR7_24_SIG,
    ADDR25      => ADDR7_25_SIG,
    ADDR26      => ADDR7_26_SIG,
    ADDR27      => ADDR7_27_SIG,
    ADDR28      => ADDR7_28_SIG,
    ADDR29      => ADDR7_29_SIG,
    ADDR30      => ADDR7_30_SIG,
    ADDR31      => ADDR7_31_SIG,
    DOUT        => VM7_OUT_SIG
);

VM8_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM8_DATA0_SIG,
    ROM1_DATA   => ROM8_DATA1_SIG,
    ROM2_DATA   => ROM8_DATA2_SIG,
    ROM3_DATA   => ROM8_DATA3_SIG,
    ROM4_DATA   => ROM8_DATA4_SIG,
    ROM5_DATA   => ROM8_DATA5_SIG,
    ROM6_DATA   => ROM8_DATA6_SIG,
    ROM7_DATA   => ROM8_DATA7_SIG,
    ROM8_DATA   => ROM8_DATA8_SIG,
    ROM9_DATA   => ROM8_DATA9_SIG,
    ROM10_DATA  => ROM8_DATA10_SIG,
    ROM11_DATA  => ROM8_DATA11_SIG,
    ROM12_DATA  => ROM8_DATA12_SIG,
    ROM13_DATA  => ROM8_DATA13_SIG,
    ROM14_DATA  => ROM8_DATA14_SIG,
    ROM15_DATA  => ROM8_DATA15_SIG,
    ROM16_DATA  => ROM8_DATA16_SIG,
    ROM17_DATA  => ROM8_DATA17_SIG,
    ROM18_DATA  => ROM8_DATA18_SIG,
    ROM19_DATA  => ROM8_DATA19_SIG,
    ROM20_DATA  => ROM8_DATA20_SIG,
    ROM21_DATA  => ROM8_DATA21_SIG,
    ROM22_DATA  => ROM8_DATA22_SIG,
    ROM23_DATA  => ROM8_DATA23_SIG,
    ROM24_DATA  => ROM8_DATA24_SIG,
    ROM25_DATA  => ROM8_DATA25_SIG,
    ROM26_DATA  => ROM8_DATA26_SIG,
    ROM27_DATA  => ROM8_DATA27_SIG,
    ROM28_DATA  => ROM8_DATA28_SIG,
    ROM29_DATA  => ROM8_DATA29_SIG,
    ROM30_DATA  => ROM8_DATA30_SIG,
    ROM31_DATA  => ROM8_DATA31_SIG,
    ADDR0       => ADDR8_0_SIG,
    ADDR1       => ADDR8_1_SIG,
    ADDR2       => ADDR8_2_SIG,
    ADDR3       => ADDR8_3_SIG,
    ADDR4       => ADDR8_4_SIG,
    ADDR5       => ADDR8_5_SIG,
    ADDR6       => ADDR8_6_SIG,
    ADDR7       => ADDR8_7_SIG,
    ADDR8       => ADDR8_8_SIG,
    ADDR9       => ADDR8_9_SIG,
    ADDR10      => ADDR8_10_SIG,
    ADDR11      => ADDR8_11_SIG,
    ADDR12      => ADDR8_12_SIG,
    ADDR13      => ADDR8_13_SIG,
    ADDR14      => ADDR8_14_SIG,
    ADDR15      => ADDR8_15_SIG,
    ADDR16      => ADDR8_16_SIG,
    ADDR17      => ADDR8_17_SIG,
    ADDR18      => ADDR8_18_SIG,
    ADDR19      => ADDR8_19_SIG,
    ADDR20      => ADDR8_20_SIG,
    ADDR21      => ADDR8_21_SIG,
    ADDR22      => ADDR8_22_SIG,
    ADDR23      => ADDR8_23_SIG,
    ADDR24      => ADDR8_24_SIG,
    ADDR25      => ADDR8_25_SIG,
    ADDR26      => ADDR8_26_SIG,
    ADDR27      => ADDR8_27_SIG,
    ADDR28      => ADDR8_28_SIG,
    ADDR29      => ADDR8_29_SIG,
    ADDR30      => ADDR8_30_SIG,
    ADDR31      => ADDR8_31_SIG,
    DOUT        => VM8_OUT_SIG
);

VM9_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM9_DATA0_SIG,
    ROM1_DATA   => ROM9_DATA1_SIG,
    ROM2_DATA   => ROM9_DATA2_SIG,
    ROM3_DATA   => ROM9_DATA3_SIG,
    ROM4_DATA   => ROM9_DATA4_SIG,
    ROM5_DATA   => ROM9_DATA5_SIG,
    ROM6_DATA   => ROM9_DATA6_SIG,
    ROM7_DATA   => ROM9_DATA7_SIG,
    ROM8_DATA   => ROM9_DATA8_SIG,
    ROM9_DATA   => ROM9_DATA9_SIG,
    ROM10_DATA  => ROM9_DATA10_SIG,
    ROM11_DATA  => ROM9_DATA11_SIG,
    ROM12_DATA  => ROM9_DATA12_SIG,
    ROM13_DATA  => ROM9_DATA13_SIG,
    ROM14_DATA  => ROM9_DATA14_SIG,
    ROM15_DATA  => ROM9_DATA15_SIG,
    ROM16_DATA  => ROM9_DATA16_SIG,
    ROM17_DATA  => ROM9_DATA17_SIG,
    ROM18_DATA  => ROM9_DATA18_SIG,
    ROM19_DATA  => ROM9_DATA19_SIG,
    ROM20_DATA  => ROM9_DATA20_SIG,
    ROM21_DATA  => ROM9_DATA21_SIG,
    ROM22_DATA  => ROM9_DATA22_SIG,
    ROM23_DATA  => ROM9_DATA23_SIG,
    ROM24_DATA  => ROM9_DATA24_SIG,
    ROM25_DATA  => ROM9_DATA25_SIG,
    ROM26_DATA  => ROM9_DATA26_SIG,
    ROM27_DATA  => ROM9_DATA27_SIG,
    ROM28_DATA  => ROM9_DATA28_SIG,
    ROM29_DATA  => ROM9_DATA29_SIG,
    ROM30_DATA  => ROM9_DATA30_SIG,
    ROM31_DATA  => ROM9_DATA31_SIG,
    ADDR0       => ADDR9_0_SIG,
    ADDR1       => ADDR9_1_SIG,
    ADDR2       => ADDR9_2_SIG,
    ADDR3       => ADDR9_3_SIG,
    ADDR4       => ADDR9_4_SIG,
    ADDR5       => ADDR9_5_SIG,
    ADDR6       => ADDR9_6_SIG,
    ADDR7       => ADDR9_7_SIG,
    ADDR8       => ADDR9_8_SIG,
    ADDR9       => ADDR9_9_SIG,
    ADDR10      => ADDR9_10_SIG,
    ADDR11      => ADDR9_11_SIG,
    ADDR12      => ADDR9_12_SIG,
    ADDR13      => ADDR9_13_SIG,
    ADDR14      => ADDR9_14_SIG,
    ADDR15      => ADDR9_15_SIG,
    ADDR16      => ADDR9_16_SIG,
    ADDR17      => ADDR9_17_SIG,
    ADDR18      => ADDR9_18_SIG,
    ADDR19      => ADDR9_19_SIG,
    ADDR20      => ADDR9_20_SIG,
    ADDR21      => ADDR9_21_SIG,
    ADDR22      => ADDR9_22_SIG,
    ADDR23      => ADDR9_23_SIG,
    ADDR24      => ADDR9_24_SIG,
    ADDR25      => ADDR9_25_SIG,
    ADDR26      => ADDR9_26_SIG,
    ADDR27      => ADDR9_27_SIG,
    ADDR28      => ADDR9_28_SIG,
    ADDR29      => ADDR9_29_SIG,
    ADDR30      => ADDR9_30_SIG,
    ADDR31      => ADDR9_31_SIG,
    DOUT        => VM9_OUT_SIG
);

VM10_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM10_DATA0_SIG,
    ROM1_DATA   => ROM10_DATA1_SIG,
    ROM2_DATA   => ROM10_DATA2_SIG,
    ROM3_DATA   => ROM10_DATA3_SIG,
    ROM4_DATA   => ROM10_DATA4_SIG,
    ROM5_DATA   => ROM10_DATA5_SIG,
    ROM6_DATA   => ROM10_DATA6_SIG,
    ROM7_DATA   => ROM10_DATA7_SIG,
    ROM8_DATA   => ROM10_DATA8_SIG,
    ROM9_DATA   => ROM10_DATA9_SIG,
    ROM10_DATA  => ROM10_DATA10_SIG,
    ROM11_DATA  => ROM10_DATA11_SIG,
    ROM12_DATA  => ROM10_DATA12_SIG,
    ROM13_DATA  => ROM10_DATA13_SIG,
    ROM14_DATA  => ROM10_DATA14_SIG,
    ROM15_DATA  => ROM10_DATA15_SIG,
    ROM16_DATA  => ROM10_DATA16_SIG,
    ROM17_DATA  => ROM10_DATA17_SIG,
    ROM18_DATA  => ROM10_DATA18_SIG,
    ROM19_DATA  => ROM10_DATA19_SIG,
    ROM20_DATA  => ROM10_DATA20_SIG,
    ROM21_DATA  => ROM10_DATA21_SIG,
    ROM22_DATA  => ROM10_DATA22_SIG,
    ROM23_DATA  => ROM10_DATA23_SIG,
    ROM24_DATA  => ROM10_DATA24_SIG,
    ROM25_DATA  => ROM10_DATA25_SIG,
    ROM26_DATA  => ROM10_DATA26_SIG,
    ROM27_DATA  => ROM10_DATA27_SIG,
    ROM28_DATA  => ROM10_DATA28_SIG,
    ROM29_DATA  => ROM10_DATA29_SIG,
    ROM30_DATA  => ROM10_DATA30_SIG,
    ROM31_DATA  => ROM10_DATA31_SIG,
    ADDR0       => ADDR10_0_SIG,
    ADDR1       => ADDR10_1_SIG,
    ADDR2       => ADDR10_2_SIG,
    ADDR3       => ADDR10_3_SIG,
    ADDR4       => ADDR10_4_SIG,
    ADDR5       => ADDR10_5_SIG,
    ADDR6       => ADDR10_6_SIG,
    ADDR7       => ADDR10_7_SIG,
    ADDR8       => ADDR10_8_SIG,
    ADDR9       => ADDR10_9_SIG,
    ADDR10      => ADDR10_10_SIG,
    ADDR11      => ADDR10_11_SIG,
    ADDR12      => ADDR10_12_SIG,
    ADDR13      => ADDR10_13_SIG,
    ADDR14      => ADDR10_14_SIG,
    ADDR15      => ADDR10_15_SIG,
    ADDR16      => ADDR10_16_SIG,
    ADDR17      => ADDR10_17_SIG,
    ADDR18      => ADDR10_18_SIG,
    ADDR19      => ADDR10_19_SIG,
    ADDR20      => ADDR10_20_SIG,
    ADDR21      => ADDR10_21_SIG,
    ADDR22      => ADDR10_22_SIG,
    ADDR23      => ADDR10_23_SIG,
    ADDR24      => ADDR10_24_SIG,
    ADDR25      => ADDR10_25_SIG,
    ADDR26      => ADDR10_26_SIG,
    ADDR27      => ADDR10_27_SIG,
    ADDR28      => ADDR10_28_SIG,
    ADDR29      => ADDR10_29_SIG,
    ADDR30      => ADDR10_30_SIG,
    ADDR31      => ADDR10_31_SIG,
    DOUT        => VM10_OUT_SIG
);

VM11_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM11_DATA0_SIG,
    ROM1_DATA   => ROM11_DATA1_SIG,
    ROM2_DATA   => ROM11_DATA2_SIG,
    ROM3_DATA   => ROM11_DATA3_SIG,
    ROM4_DATA   => ROM11_DATA4_SIG,
    ROM5_DATA   => ROM11_DATA5_SIG,
    ROM6_DATA   => ROM11_DATA6_SIG,
    ROM7_DATA   => ROM11_DATA7_SIG,
    ROM8_DATA   => ROM11_DATA8_SIG,
    ROM9_DATA   => ROM11_DATA9_SIG,
    ROM10_DATA  => ROM11_DATA10_SIG,
    ROM11_DATA  => ROM11_DATA11_SIG,
    ROM12_DATA  => ROM11_DATA12_SIG,
    ROM13_DATA  => ROM11_DATA13_SIG,
    ROM14_DATA  => ROM11_DATA14_SIG,
    ROM15_DATA  => ROM11_DATA15_SIG,
    ROM16_DATA  => ROM11_DATA16_SIG,
    ROM17_DATA  => ROM11_DATA17_SIG,
    ROM18_DATA  => ROM11_DATA18_SIG,
    ROM19_DATA  => ROM11_DATA19_SIG,
    ROM20_DATA  => ROM11_DATA20_SIG,
    ROM21_DATA  => ROM11_DATA21_SIG,
    ROM22_DATA  => ROM11_DATA22_SIG,
    ROM23_DATA  => ROM11_DATA23_SIG,
    ROM24_DATA  => ROM11_DATA24_SIG,
    ROM25_DATA  => ROM11_DATA25_SIG,
    ROM26_DATA  => ROM11_DATA26_SIG,
    ROM27_DATA  => ROM11_DATA27_SIG,
    ROM28_DATA  => ROM11_DATA28_SIG,
    ROM29_DATA  => ROM11_DATA29_SIG,
    ROM30_DATA  => ROM11_DATA30_SIG,
    ROM31_DATA  => ROM11_DATA31_SIG,
    ADDR0       => ADDR11_0_SIG,
    ADDR1       => ADDR11_1_SIG,
    ADDR2       => ADDR11_2_SIG,
    ADDR3       => ADDR11_3_SIG,
    ADDR4       => ADDR11_4_SIG,
    ADDR5       => ADDR11_5_SIG,
    ADDR6       => ADDR11_6_SIG,
    ADDR7       => ADDR11_7_SIG,
    ADDR8       => ADDR11_8_SIG,
    ADDR9       => ADDR11_9_SIG,
    ADDR10      => ADDR11_10_SIG,
    ADDR11      => ADDR11_11_SIG,
    ADDR12      => ADDR11_12_SIG,
    ADDR13      => ADDR11_13_SIG,
    ADDR14      => ADDR11_14_SIG,
    ADDR15      => ADDR11_15_SIG,
    ADDR16      => ADDR11_16_SIG,
    ADDR17      => ADDR11_17_SIG,
    ADDR18      => ADDR11_18_SIG,
    ADDR19      => ADDR11_19_SIG,
    ADDR20      => ADDR11_20_SIG,
    ADDR21      => ADDR11_21_SIG,
    ADDR22      => ADDR11_22_SIG,
    ADDR23      => ADDR11_23_SIG,
    ADDR24      => ADDR11_24_SIG,
    ADDR25      => ADDR11_25_SIG,
    ADDR26      => ADDR11_26_SIG,
    ADDR27      => ADDR11_27_SIG,
    ADDR28      => ADDR11_28_SIG,
    ADDR29      => ADDR11_29_SIG,
    ADDR30      => ADDR11_30_SIG,
    ADDR31      => ADDR11_31_SIG,
    DOUT        => VM11_OUT_SIG
);

VM12_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM12_DATA0_SIG,
    ROM1_DATA   => ROM12_DATA1_SIG,
    ROM2_DATA   => ROM12_DATA2_SIG,
    ROM3_DATA   => ROM12_DATA3_SIG,
    ROM4_DATA   => ROM12_DATA4_SIG,
    ROM5_DATA   => ROM12_DATA5_SIG,
    ROM6_DATA   => ROM12_DATA6_SIG,
    ROM7_DATA   => ROM12_DATA7_SIG,
    ROM8_DATA   => ROM12_DATA8_SIG,
    ROM9_DATA   => ROM12_DATA9_SIG,
    ROM10_DATA  => ROM12_DATA10_SIG,
    ROM11_DATA  => ROM12_DATA11_SIG,
    ROM12_DATA  => ROM12_DATA12_SIG,
    ROM13_DATA  => ROM12_DATA13_SIG,
    ROM14_DATA  => ROM12_DATA14_SIG,
    ROM15_DATA  => ROM12_DATA15_SIG,
    ROM16_DATA  => ROM12_DATA16_SIG,
    ROM17_DATA  => ROM12_DATA17_SIG,
    ROM18_DATA  => ROM12_DATA18_SIG,
    ROM19_DATA  => ROM12_DATA19_SIG,
    ROM20_DATA  => ROM12_DATA20_SIG,
    ROM21_DATA  => ROM12_DATA21_SIG,
    ROM22_DATA  => ROM12_DATA22_SIG,
    ROM23_DATA  => ROM12_DATA23_SIG,
    ROM24_DATA  => ROM12_DATA24_SIG,
    ROM25_DATA  => ROM12_DATA25_SIG,
    ROM26_DATA  => ROM12_DATA26_SIG,
    ROM27_DATA  => ROM12_DATA27_SIG,
    ROM28_DATA  => ROM12_DATA28_SIG,
    ROM29_DATA  => ROM12_DATA29_SIG,
    ROM30_DATA  => ROM12_DATA30_SIG,
    ROM31_DATA  => ROM12_DATA31_SIG,
    ADDR0       => ADDR12_0_SIG,
    ADDR1       => ADDR12_1_SIG,
    ADDR2       => ADDR12_2_SIG,
    ADDR3       => ADDR12_3_SIG,
    ADDR4       => ADDR12_4_SIG,
    ADDR5       => ADDR12_5_SIG,
    ADDR6       => ADDR12_6_SIG,
    ADDR7       => ADDR12_7_SIG,
    ADDR8       => ADDR12_8_SIG,
    ADDR9       => ADDR12_9_SIG,
    ADDR10      => ADDR12_10_SIG,
    ADDR11      => ADDR12_11_SIG,
    ADDR12      => ADDR12_12_SIG,
    ADDR13      => ADDR12_13_SIG,
    ADDR14      => ADDR12_14_SIG,
    ADDR15      => ADDR12_15_SIG,
    ADDR16      => ADDR12_16_SIG,
    ADDR17      => ADDR12_17_SIG,
    ADDR18      => ADDR12_18_SIG,
    ADDR19      => ADDR12_19_SIG,
    ADDR20      => ADDR12_20_SIG,
    ADDR21      => ADDR12_21_SIG,
    ADDR22      => ADDR12_22_SIG,
    ADDR23      => ADDR12_23_SIG,
    ADDR24      => ADDR12_24_SIG,
    ADDR25      => ADDR12_25_SIG,
    ADDR26      => ADDR12_26_SIG,
    ADDR27      => ADDR12_27_SIG,
    ADDR28      => ADDR12_28_SIG,
    ADDR29      => ADDR12_29_SIG,
    ADDR30      => ADDR12_30_SIG,
    ADDR31      => ADDR12_31_SIG,
    DOUT        => VM12_OUT_SIG
);

VM13_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM13_DATA0_SIG,
    ROM1_DATA   => ROM13_DATA1_SIG,
    ROM2_DATA   => ROM13_DATA2_SIG,
    ROM3_DATA   => ROM13_DATA3_SIG,
    ROM4_DATA   => ROM13_DATA4_SIG,
    ROM5_DATA   => ROM13_DATA5_SIG,
    ROM6_DATA   => ROM13_DATA6_SIG,
    ROM7_DATA   => ROM13_DATA7_SIG,
    ROM8_DATA   => ROM13_DATA8_SIG,
    ROM9_DATA   => ROM13_DATA9_SIG,
    ROM10_DATA  => ROM13_DATA10_SIG,
    ROM11_DATA  => ROM13_DATA11_SIG,
    ROM12_DATA  => ROM13_DATA12_SIG,
    ROM13_DATA  => ROM13_DATA13_SIG,
    ROM14_DATA  => ROM13_DATA14_SIG,
    ROM15_DATA  => ROM13_DATA15_SIG,
    ROM16_DATA  => ROM13_DATA16_SIG,
    ROM17_DATA  => ROM13_DATA17_SIG,
    ROM18_DATA  => ROM13_DATA18_SIG,
    ROM19_DATA  => ROM13_DATA19_SIG,
    ROM20_DATA  => ROM13_DATA20_SIG,
    ROM21_DATA  => ROM13_DATA21_SIG,
    ROM22_DATA  => ROM13_DATA22_SIG,
    ROM23_DATA  => ROM13_DATA23_SIG,
    ROM24_DATA  => ROM13_DATA24_SIG,
    ROM25_DATA  => ROM13_DATA25_SIG,
    ROM26_DATA  => ROM13_DATA26_SIG,
    ROM27_DATA  => ROM13_DATA27_SIG,
    ROM28_DATA  => ROM13_DATA28_SIG,
    ROM29_DATA  => ROM13_DATA29_SIG,
    ROM30_DATA  => ROM13_DATA30_SIG,
    ROM31_DATA  => ROM13_DATA31_SIG,
    ADDR0       => ADDR13_0_SIG,
    ADDR1       => ADDR13_1_SIG,
    ADDR2       => ADDR13_2_SIG,
    ADDR3       => ADDR13_3_SIG,
    ADDR4       => ADDR13_4_SIG,
    ADDR5       => ADDR13_5_SIG,
    ADDR6       => ADDR13_6_SIG,
    ADDR7       => ADDR13_7_SIG,
    ADDR8       => ADDR13_8_SIG,
    ADDR9       => ADDR13_9_SIG,
    ADDR10      => ADDR13_10_SIG,
    ADDR11      => ADDR13_11_SIG,
    ADDR12      => ADDR13_12_SIG,
    ADDR13      => ADDR13_13_SIG,
    ADDR14      => ADDR13_14_SIG,
    ADDR15      => ADDR13_15_SIG,
    ADDR16      => ADDR13_16_SIG,
    ADDR17      => ADDR13_17_SIG,
    ADDR18      => ADDR13_18_SIG,
    ADDR19      => ADDR13_19_SIG,
    ADDR20      => ADDR13_20_SIG,
    ADDR21      => ADDR13_21_SIG,
    ADDR22      => ADDR13_22_SIG,
    ADDR23      => ADDR13_23_SIG,
    ADDR24      => ADDR13_24_SIG,
    ADDR25      => ADDR13_25_SIG,
    ADDR26      => ADDR13_26_SIG,
    ADDR27      => ADDR13_27_SIG,
    ADDR28      => ADDR13_28_SIG,
    ADDR29      => ADDR13_29_SIG,
    ADDR30      => ADDR13_30_SIG,
    ADDR31      => ADDR13_31_SIG,
    DOUT        => VM13_OUT_SIG
);

VM14_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM14_DATA0_SIG,
    ROM1_DATA   => ROM14_DATA1_SIG,
    ROM2_DATA   => ROM14_DATA2_SIG,
    ROM3_DATA   => ROM14_DATA3_SIG,
    ROM4_DATA   => ROM14_DATA4_SIG,
    ROM5_DATA   => ROM14_DATA5_SIG,
    ROM6_DATA   => ROM14_DATA6_SIG,
    ROM7_DATA   => ROM14_DATA7_SIG,
    ROM8_DATA   => ROM14_DATA8_SIG,
    ROM9_DATA   => ROM14_DATA9_SIG,
    ROM10_DATA  => ROM14_DATA10_SIG,
    ROM11_DATA  => ROM14_DATA11_SIG,
    ROM12_DATA  => ROM14_DATA12_SIG,
    ROM13_DATA  => ROM14_DATA13_SIG,
    ROM14_DATA  => ROM14_DATA14_SIG,
    ROM15_DATA  => ROM14_DATA15_SIG,
    ROM16_DATA  => ROM14_DATA16_SIG,
    ROM17_DATA  => ROM14_DATA17_SIG,
    ROM18_DATA  => ROM14_DATA18_SIG,
    ROM19_DATA  => ROM14_DATA19_SIG,
    ROM20_DATA  => ROM14_DATA20_SIG,
    ROM21_DATA  => ROM14_DATA21_SIG,
    ROM22_DATA  => ROM14_DATA22_SIG,
    ROM23_DATA  => ROM14_DATA23_SIG,
    ROM24_DATA  => ROM14_DATA24_SIG,
    ROM25_DATA  => ROM14_DATA25_SIG,
    ROM26_DATA  => ROM14_DATA26_SIG,
    ROM27_DATA  => ROM14_DATA27_SIG,
    ROM28_DATA  => ROM14_DATA28_SIG,
    ROM29_DATA  => ROM14_DATA29_SIG,
    ROM30_DATA  => ROM14_DATA30_SIG,
    ROM31_DATA  => ROM14_DATA31_SIG,
    ADDR0       => ADDR14_0_SIG,
    ADDR1       => ADDR14_1_SIG,
    ADDR2       => ADDR14_2_SIG,
    ADDR3       => ADDR14_3_SIG,
    ADDR4       => ADDR14_4_SIG,
    ADDR5       => ADDR14_5_SIG,
    ADDR6       => ADDR14_6_SIG,
    ADDR7       => ADDR14_7_SIG,
    ADDR8       => ADDR14_8_SIG,
    ADDR9       => ADDR14_9_SIG,
    ADDR10      => ADDR14_10_SIG,
    ADDR11      => ADDR14_11_SIG,
    ADDR12      => ADDR14_12_SIG,
    ADDR13      => ADDR14_13_SIG,
    ADDR14      => ADDR14_14_SIG,
    ADDR15      => ADDR14_15_SIG,
    ADDR16      => ADDR14_16_SIG,
    ADDR17      => ADDR14_17_SIG,
    ADDR18      => ADDR14_18_SIG,
    ADDR19      => ADDR14_19_SIG,
    ADDR20      => ADDR14_20_SIG,
    ADDR21      => ADDR14_21_SIG,
    ADDR22      => ADDR14_22_SIG,
    ADDR23      => ADDR14_23_SIG,
    ADDR24      => ADDR14_24_SIG,
    ADDR25      => ADDR14_25_SIG,
    ADDR26      => ADDR14_26_SIG,
    ADDR27      => ADDR14_27_SIG,
    ADDR28      => ADDR14_28_SIG,
    ADDR29      => ADDR14_29_SIG,
    ADDR30      => ADDR14_30_SIG,
    ADDR31      => ADDR14_31_SIG,
    DOUT        => VM14_OUT_SIG
);

VM15_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM15_DATA0_SIG,
    ROM1_DATA   => ROM15_DATA1_SIG,
    ROM2_DATA   => ROM15_DATA2_SIG,
    ROM3_DATA   => ROM15_DATA3_SIG,
    ROM4_DATA   => ROM15_DATA4_SIG,
    ROM5_DATA   => ROM15_DATA5_SIG,
    ROM6_DATA   => ROM15_DATA6_SIG,
    ROM7_DATA   => ROM15_DATA7_SIG,
    ROM8_DATA   => ROM15_DATA8_SIG,
    ROM9_DATA   => ROM15_DATA9_SIG,
    ROM10_DATA  => ROM15_DATA10_SIG,
    ROM11_DATA  => ROM15_DATA11_SIG,
    ROM12_DATA  => ROM15_DATA12_SIG,
    ROM13_DATA  => ROM15_DATA13_SIG,
    ROM14_DATA  => ROM15_DATA14_SIG,
    ROM15_DATA  => ROM15_DATA15_SIG,
    ROM16_DATA  => ROM15_DATA16_SIG,
    ROM17_DATA  => ROM15_DATA17_SIG,
    ROM18_DATA  => ROM15_DATA18_SIG,
    ROM19_DATA  => ROM15_DATA19_SIG,
    ROM20_DATA  => ROM15_DATA20_SIG,
    ROM21_DATA  => ROM15_DATA21_SIG,
    ROM22_DATA  => ROM15_DATA22_SIG,
    ROM23_DATA  => ROM15_DATA23_SIG,
    ROM24_DATA  => ROM15_DATA24_SIG,
    ROM25_DATA  => ROM15_DATA25_SIG,
    ROM26_DATA  => ROM15_DATA26_SIG,
    ROM27_DATA  => ROM15_DATA27_SIG,
    ROM28_DATA  => ROM15_DATA28_SIG,
    ROM29_DATA  => ROM15_DATA29_SIG,
    ROM30_DATA  => ROM15_DATA30_SIG,
    ROM31_DATA  => ROM15_DATA31_SIG,
    ADDR0       => ADDR15_0_SIG,
    ADDR1       => ADDR15_1_SIG,
    ADDR2       => ADDR15_2_SIG,
    ADDR3       => ADDR15_3_SIG,
    ADDR4       => ADDR15_4_SIG,
    ADDR5       => ADDR15_5_SIG,
    ADDR6       => ADDR15_6_SIG,
    ADDR7       => ADDR15_7_SIG,
    ADDR8       => ADDR15_8_SIG,
    ADDR9       => ADDR15_9_SIG,
    ADDR10      => ADDR15_10_SIG,
    ADDR11      => ADDR15_11_SIG,
    ADDR12      => ADDR15_12_SIG,
    ADDR13      => ADDR15_13_SIG,
    ADDR14      => ADDR15_14_SIG,
    ADDR15      => ADDR15_15_SIG,
    ADDR16      => ADDR15_16_SIG,
    ADDR17      => ADDR15_17_SIG,
    ADDR18      => ADDR15_18_SIG,
    ADDR19      => ADDR15_19_SIG,
    ADDR20      => ADDR15_20_SIG,
    ADDR21      => ADDR15_21_SIG,
    ADDR22      => ADDR15_22_SIG,
    ADDR23      => ADDR15_23_SIG,
    ADDR24      => ADDR15_24_SIG,
    ADDR25      => ADDR15_25_SIG,
    ADDR26      => ADDR15_26_SIG,
    ADDR27      => ADDR15_27_SIG,
    ADDR28      => ADDR15_28_SIG,
    ADDR29      => ADDR15_29_SIG,
    ADDR30      => ADDR15_30_SIG,
    ADDR31      => ADDR15_31_SIG,
    DOUT        => VM15_OUT_SIG
);

VM16_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM16_DATA0_SIG,
    ROM1_DATA   => ROM16_DATA1_SIG,
    ROM2_DATA   => ROM16_DATA2_SIG,
    ROM3_DATA   => ROM16_DATA3_SIG,
    ROM4_DATA   => ROM16_DATA4_SIG,
    ROM5_DATA   => ROM16_DATA5_SIG,
    ROM6_DATA   => ROM16_DATA6_SIG,
    ROM7_DATA   => ROM16_DATA7_SIG,
    ROM8_DATA   => ROM16_DATA8_SIG,
    ROM9_DATA   => ROM16_DATA9_SIG,
    ROM10_DATA  => ROM16_DATA10_SIG,
    ROM11_DATA  => ROM16_DATA11_SIG,
    ROM12_DATA  => ROM16_DATA12_SIG,
    ROM13_DATA  => ROM16_DATA13_SIG,
    ROM14_DATA  => ROM16_DATA14_SIG,
    ROM15_DATA  => ROM16_DATA15_SIG,
    ROM16_DATA  => ROM16_DATA16_SIG,
    ROM17_DATA  => ROM16_DATA17_SIG,
    ROM18_DATA  => ROM16_DATA18_SIG,
    ROM19_DATA  => ROM16_DATA19_SIG,
    ROM20_DATA  => ROM16_DATA20_SIG,
    ROM21_DATA  => ROM16_DATA21_SIG,
    ROM22_DATA  => ROM16_DATA22_SIG,
    ROM23_DATA  => ROM16_DATA23_SIG,
    ROM24_DATA  => ROM16_DATA24_SIG,
    ROM25_DATA  => ROM16_DATA25_SIG,
    ROM26_DATA  => ROM16_DATA26_SIG,
    ROM27_DATA  => ROM16_DATA27_SIG,
    ROM28_DATA  => ROM16_DATA28_SIG,
    ROM29_DATA  => ROM16_DATA29_SIG,
    ROM30_DATA  => ROM16_DATA30_SIG,
    ROM31_DATA  => ROM16_DATA31_SIG,
    ADDR0       => ADDR16_0_SIG,
    ADDR1       => ADDR16_1_SIG,
    ADDR2       => ADDR16_2_SIG,
    ADDR3       => ADDR16_3_SIG,
    ADDR4       => ADDR16_4_SIG,
    ADDR5       => ADDR16_5_SIG,
    ADDR6       => ADDR16_6_SIG,
    ADDR7       => ADDR16_7_SIG,
    ADDR8       => ADDR16_8_SIG,
    ADDR9       => ADDR16_9_SIG,
    ADDR10      => ADDR16_10_SIG,
    ADDR11      => ADDR16_11_SIG,
    ADDR12      => ADDR16_12_SIG,
    ADDR13      => ADDR16_13_SIG,
    ADDR14      => ADDR16_14_SIG,
    ADDR15      => ADDR16_15_SIG,
    ADDR16      => ADDR16_16_SIG,
    ADDR17      => ADDR16_17_SIG,
    ADDR18      => ADDR16_18_SIG,
    ADDR19      => ADDR16_19_SIG,
    ADDR20      => ADDR16_20_SIG,
    ADDR21      => ADDR16_21_SIG,
    ADDR22      => ADDR16_22_SIG,
    ADDR23      => ADDR16_23_SIG,
    ADDR24      => ADDR16_24_SIG,
    ADDR25      => ADDR16_25_SIG,
    ADDR26      => ADDR16_26_SIG,
    ADDR27      => ADDR16_27_SIG,
    ADDR28      => ADDR16_28_SIG,
    ADDR29      => ADDR16_29_SIG,
    ADDR30      => ADDR16_30_SIG,
    ADDR31      => ADDR16_31_SIG,
    DOUT        => VM16_OUT_SIG
);

VM17_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM17_DATA0_SIG,
    ROM1_DATA   => ROM17_DATA1_SIG,
    ROM2_DATA   => ROM17_DATA2_SIG,
    ROM3_DATA   => ROM17_DATA3_SIG,
    ROM4_DATA   => ROM17_DATA4_SIG,
    ROM5_DATA   => ROM17_DATA5_SIG,
    ROM6_DATA   => ROM17_DATA6_SIG,
    ROM7_DATA   => ROM17_DATA7_SIG,
    ROM8_DATA   => ROM17_DATA8_SIG,
    ROM9_DATA   => ROM17_DATA9_SIG,
    ROM10_DATA  => ROM17_DATA10_SIG,
    ROM11_DATA  => ROM17_DATA11_SIG,
    ROM12_DATA  => ROM17_DATA12_SIG,
    ROM13_DATA  => ROM17_DATA13_SIG,
    ROM14_DATA  => ROM17_DATA14_SIG,
    ROM15_DATA  => ROM17_DATA15_SIG,
    ROM16_DATA  => ROM17_DATA16_SIG,
    ROM17_DATA  => ROM17_DATA17_SIG,
    ROM18_DATA  => ROM17_DATA18_SIG,
    ROM19_DATA  => ROM17_DATA19_SIG,
    ROM20_DATA  => ROM17_DATA20_SIG,
    ROM21_DATA  => ROM17_DATA21_SIG,
    ROM22_DATA  => ROM17_DATA22_SIG,
    ROM23_DATA  => ROM17_DATA23_SIG,
    ROM24_DATA  => ROM17_DATA24_SIG,
    ROM25_DATA  => ROM17_DATA25_SIG,
    ROM26_DATA  => ROM17_DATA26_SIG,
    ROM27_DATA  => ROM17_DATA27_SIG,
    ROM28_DATA  => ROM17_DATA28_SIG,
    ROM29_DATA  => ROM17_DATA29_SIG,
    ROM30_DATA  => ROM17_DATA30_SIG,
    ROM31_DATA  => ROM17_DATA31_SIG,
    ADDR0       => ADDR17_0_SIG,
    ADDR1       => ADDR17_1_SIG,
    ADDR2       => ADDR17_2_SIG,
    ADDR3       => ADDR17_3_SIG,
    ADDR4       => ADDR17_4_SIG,
    ADDR5       => ADDR17_5_SIG,
    ADDR6       => ADDR17_6_SIG,
    ADDR7       => ADDR17_7_SIG,
    ADDR8       => ADDR17_8_SIG,
    ADDR9       => ADDR17_9_SIG,
    ADDR10      => ADDR17_10_SIG,
    ADDR11      => ADDR17_11_SIG,
    ADDR12      => ADDR17_12_SIG,
    ADDR13      => ADDR17_13_SIG,
    ADDR14      => ADDR17_14_SIG,
    ADDR15      => ADDR17_15_SIG,
    ADDR16      => ADDR17_16_SIG,
    ADDR17      => ADDR17_17_SIG,
    ADDR18      => ADDR17_18_SIG,
    ADDR19      => ADDR17_19_SIG,
    ADDR20      => ADDR17_20_SIG,
    ADDR21      => ADDR17_21_SIG,
    ADDR22      => ADDR17_22_SIG,
    ADDR23      => ADDR17_23_SIG,
    ADDR24      => ADDR17_24_SIG,
    ADDR25      => ADDR17_25_SIG,
    ADDR26      => ADDR17_26_SIG,
    ADDR27      => ADDR17_27_SIG,
    ADDR28      => ADDR17_28_SIG,
    ADDR29      => ADDR17_29_SIG,
    ADDR30      => ADDR17_30_SIG,
    ADDR31      => ADDR17_31_SIG,
    DOUT        => VM17_OUT_SIG
);

VM18_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM18_DATA0_SIG,
    ROM1_DATA   => ROM18_DATA1_SIG,
    ROM2_DATA   => ROM18_DATA2_SIG,
    ROM3_DATA   => ROM18_DATA3_SIG,
    ROM4_DATA   => ROM18_DATA4_SIG,
    ROM5_DATA   => ROM18_DATA5_SIG,
    ROM6_DATA   => ROM18_DATA6_SIG,
    ROM7_DATA   => ROM18_DATA7_SIG,
    ROM8_DATA   => ROM18_DATA8_SIG,
    ROM9_DATA   => ROM18_DATA9_SIG,
    ROM10_DATA  => ROM18_DATA10_SIG,
    ROM11_DATA  => ROM18_DATA11_SIG,
    ROM12_DATA  => ROM18_DATA12_SIG,
    ROM13_DATA  => ROM18_DATA13_SIG,
    ROM14_DATA  => ROM18_DATA14_SIG,
    ROM15_DATA  => ROM18_DATA15_SIG,
    ROM16_DATA  => ROM18_DATA16_SIG,
    ROM17_DATA  => ROM18_DATA17_SIG,
    ROM18_DATA  => ROM18_DATA18_SIG,
    ROM19_DATA  => ROM18_DATA19_SIG,
    ROM20_DATA  => ROM18_DATA20_SIG,
    ROM21_DATA  => ROM18_DATA21_SIG,
    ROM22_DATA  => ROM18_DATA22_SIG,
    ROM23_DATA  => ROM18_DATA23_SIG,
    ROM24_DATA  => ROM18_DATA24_SIG,
    ROM25_DATA  => ROM18_DATA25_SIG,
    ROM26_DATA  => ROM18_DATA26_SIG,
    ROM27_DATA  => ROM18_DATA27_SIG,
    ROM28_DATA  => ROM18_DATA28_SIG,
    ROM29_DATA  => ROM18_DATA29_SIG,
    ROM30_DATA  => ROM18_DATA30_SIG,
    ROM31_DATA  => ROM18_DATA31_SIG,
    ADDR0       => ADDR18_0_SIG,
    ADDR1       => ADDR18_1_SIG,
    ADDR2       => ADDR18_2_SIG,
    ADDR3       => ADDR18_3_SIG,
    ADDR4       => ADDR18_4_SIG,
    ADDR5       => ADDR18_5_SIG,
    ADDR6       => ADDR18_6_SIG,
    ADDR7       => ADDR18_7_SIG,
    ADDR8       => ADDR18_8_SIG,
    ADDR9       => ADDR18_9_SIG,
    ADDR10      => ADDR18_10_SIG,
    ADDR11      => ADDR18_11_SIG,
    ADDR12      => ADDR18_12_SIG,
    ADDR13      => ADDR18_13_SIG,
    ADDR14      => ADDR18_14_SIG,
    ADDR15      => ADDR18_15_SIG,
    ADDR16      => ADDR18_16_SIG,
    ADDR17      => ADDR18_17_SIG,
    ADDR18      => ADDR18_18_SIG,
    ADDR19      => ADDR18_19_SIG,
    ADDR20      => ADDR18_20_SIG,
    ADDR21      => ADDR18_21_SIG,
    ADDR22      => ADDR18_22_SIG,
    ADDR23      => ADDR18_23_SIG,
    ADDR24      => ADDR18_24_SIG,
    ADDR25      => ADDR18_25_SIG,
    ADDR26      => ADDR18_26_SIG,
    ADDR27      => ADDR18_27_SIG,
    ADDR28      => ADDR18_28_SIG,
    ADDR29      => ADDR18_29_SIG,
    ADDR30      => ADDR18_30_SIG,
    ADDR31      => ADDR18_31_SIG,
    DOUT        => VM18_OUT_SIG
);

VM19_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM19_DATA0_SIG,
    ROM1_DATA   => ROM19_DATA1_SIG,
    ROM2_DATA   => ROM19_DATA2_SIG,
    ROM3_DATA   => ROM19_DATA3_SIG,
    ROM4_DATA   => ROM19_DATA4_SIG,
    ROM5_DATA   => ROM19_DATA5_SIG,
    ROM6_DATA   => ROM19_DATA6_SIG,
    ROM7_DATA   => ROM19_DATA7_SIG,
    ROM8_DATA   => ROM19_DATA8_SIG,
    ROM9_DATA   => ROM19_DATA9_SIG,
    ROM10_DATA  => ROM19_DATA10_SIG,
    ROM11_DATA  => ROM19_DATA11_SIG,
    ROM12_DATA  => ROM19_DATA12_SIG,
    ROM13_DATA  => ROM19_DATA13_SIG,
    ROM14_DATA  => ROM19_DATA14_SIG,
    ROM15_DATA  => ROM19_DATA15_SIG,
    ROM16_DATA  => ROM19_DATA16_SIG,
    ROM17_DATA  => ROM19_DATA17_SIG,
    ROM18_DATA  => ROM19_DATA18_SIG,
    ROM19_DATA  => ROM19_DATA19_SIG,
    ROM20_DATA  => ROM19_DATA20_SIG,
    ROM21_DATA  => ROM19_DATA21_SIG,
    ROM22_DATA  => ROM19_DATA22_SIG,
    ROM23_DATA  => ROM19_DATA23_SIG,
    ROM24_DATA  => ROM19_DATA24_SIG,
    ROM25_DATA  => ROM19_DATA25_SIG,
    ROM26_DATA  => ROM19_DATA26_SIG,
    ROM27_DATA  => ROM19_DATA27_SIG,
    ROM28_DATA  => ROM19_DATA28_SIG,
    ROM29_DATA  => ROM19_DATA29_SIG,
    ROM30_DATA  => ROM19_DATA30_SIG,
    ROM31_DATA  => ROM19_DATA31_SIG,
    ADDR0       => ADDR19_0_SIG,
    ADDR1       => ADDR19_1_SIG,
    ADDR2       => ADDR19_2_SIG,
    ADDR3       => ADDR19_3_SIG,
    ADDR4       => ADDR19_4_SIG,
    ADDR5       => ADDR19_5_SIG,
    ADDR6       => ADDR19_6_SIG,
    ADDR7       => ADDR19_7_SIG,
    ADDR8       => ADDR19_8_SIG,
    ADDR9       => ADDR19_9_SIG,
    ADDR10      => ADDR19_10_SIG,
    ADDR11      => ADDR19_11_SIG,
    ADDR12      => ADDR19_12_SIG,
    ADDR13      => ADDR19_13_SIG,
    ADDR14      => ADDR19_14_SIG,
    ADDR15      => ADDR19_15_SIG,
    ADDR16      => ADDR19_16_SIG,
    ADDR17      => ADDR19_17_SIG,
    ADDR18      => ADDR19_18_SIG,
    ADDR19      => ADDR19_19_SIG,
    ADDR20      => ADDR19_20_SIG,
    ADDR21      => ADDR19_21_SIG,
    ADDR22      => ADDR19_22_SIG,
    ADDR23      => ADDR19_23_SIG,
    ADDR24      => ADDR19_24_SIG,
    ADDR25      => ADDR19_25_SIG,
    ADDR26      => ADDR19_26_SIG,
    ADDR27      => ADDR19_27_SIG,
    ADDR28      => ADDR19_28_SIG,
    ADDR29      => ADDR19_29_SIG,
    ADDR30      => ADDR19_30_SIG,
    ADDR31      => ADDR19_31_SIG,
    DOUT        => VM19_OUT_SIG
);

VM20_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM20_DATA0_SIG,
    ROM1_DATA   => ROM20_DATA1_SIG,
    ROM2_DATA   => ROM20_DATA2_SIG,
    ROM3_DATA   => ROM20_DATA3_SIG,
    ROM4_DATA   => ROM20_DATA4_SIG,
    ROM5_DATA   => ROM20_DATA5_SIG,
    ROM6_DATA   => ROM20_DATA6_SIG,
    ROM7_DATA   => ROM20_DATA7_SIG,
    ROM8_DATA   => ROM20_DATA8_SIG,
    ROM9_DATA   => ROM20_DATA9_SIG,
    ROM10_DATA  => ROM20_DATA10_SIG,
    ROM11_DATA  => ROM20_DATA11_SIG,
    ROM12_DATA  => ROM20_DATA12_SIG,
    ROM13_DATA  => ROM20_DATA13_SIG,
    ROM14_DATA  => ROM20_DATA14_SIG,
    ROM15_DATA  => ROM20_DATA15_SIG,
    ROM16_DATA  => ROM20_DATA16_SIG,
    ROM17_DATA  => ROM20_DATA17_SIG,
    ROM18_DATA  => ROM20_DATA18_SIG,
    ROM19_DATA  => ROM20_DATA19_SIG,
    ROM20_DATA  => ROM20_DATA20_SIG,
    ROM21_DATA  => ROM20_DATA21_SIG,
    ROM22_DATA  => ROM20_DATA22_SIG,
    ROM23_DATA  => ROM20_DATA23_SIG,
    ROM24_DATA  => ROM20_DATA24_SIG,
    ROM25_DATA  => ROM20_DATA25_SIG,
    ROM26_DATA  => ROM20_DATA26_SIG,
    ROM27_DATA  => ROM20_DATA27_SIG,
    ROM28_DATA  => ROM20_DATA28_SIG,
    ROM29_DATA  => ROM20_DATA29_SIG,
    ROM30_DATA  => ROM20_DATA30_SIG,
    ROM31_DATA  => ROM20_DATA31_SIG,
    ADDR0       => ADDR20_0_SIG,
    ADDR1       => ADDR20_1_SIG,
    ADDR2       => ADDR20_2_SIG,
    ADDR3       => ADDR20_3_SIG,
    ADDR4       => ADDR20_4_SIG,
    ADDR5       => ADDR20_5_SIG,
    ADDR6       => ADDR20_6_SIG,
    ADDR7       => ADDR20_7_SIG,
    ADDR8       => ADDR20_8_SIG,
    ADDR9       => ADDR20_9_SIG,
    ADDR10      => ADDR20_10_SIG,
    ADDR11      => ADDR20_11_SIG,
    ADDR12      => ADDR20_12_SIG,
    ADDR13      => ADDR20_13_SIG,
    ADDR14      => ADDR20_14_SIG,
    ADDR15      => ADDR20_15_SIG,
    ADDR16      => ADDR20_16_SIG,
    ADDR17      => ADDR20_17_SIG,
    ADDR18      => ADDR20_18_SIG,
    ADDR19      => ADDR20_19_SIG,
    ADDR20      => ADDR20_20_SIG,
    ADDR21      => ADDR20_21_SIG,
    ADDR22      => ADDR20_22_SIG,
    ADDR23      => ADDR20_23_SIG,
    ADDR24      => ADDR20_24_SIG,
    ADDR25      => ADDR20_25_SIG,
    ADDR26      => ADDR20_26_SIG,
    ADDR27      => ADDR20_27_SIG,
    ADDR28      => ADDR20_28_SIG,
    ADDR29      => ADDR20_29_SIG,
    ADDR30      => ADDR20_30_SIG,
    ADDR31      => ADDR20_31_SIG,
    DOUT        => VM20_OUT_SIG
);

VM21_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM21_DATA0_SIG,
    ROM1_DATA   => ROM21_DATA1_SIG,
    ROM2_DATA   => ROM21_DATA2_SIG,
    ROM3_DATA   => ROM21_DATA3_SIG,
    ROM4_DATA   => ROM21_DATA4_SIG,
    ROM5_DATA   => ROM21_DATA5_SIG,
    ROM6_DATA   => ROM21_DATA6_SIG,
    ROM7_DATA   => ROM21_DATA7_SIG,
    ROM8_DATA   => ROM21_DATA8_SIG,
    ROM9_DATA   => ROM21_DATA9_SIG,
    ROM10_DATA  => ROM21_DATA10_SIG,
    ROM11_DATA  => ROM21_DATA11_SIG,
    ROM12_DATA  => ROM21_DATA12_SIG,
    ROM13_DATA  => ROM21_DATA13_SIG,
    ROM14_DATA  => ROM21_DATA14_SIG,
    ROM15_DATA  => ROM21_DATA15_SIG,
    ROM16_DATA  => ROM21_DATA16_SIG,
    ROM17_DATA  => ROM21_DATA17_SIG,
    ROM18_DATA  => ROM21_DATA18_SIG,
    ROM19_DATA  => ROM21_DATA19_SIG,
    ROM20_DATA  => ROM21_DATA20_SIG,
    ROM21_DATA  => ROM21_DATA21_SIG,
    ROM22_DATA  => ROM21_DATA22_SIG,
    ROM23_DATA  => ROM21_DATA23_SIG,
    ROM24_DATA  => ROM21_DATA24_SIG,
    ROM25_DATA  => ROM21_DATA25_SIG,
    ROM26_DATA  => ROM21_DATA26_SIG,
    ROM27_DATA  => ROM21_DATA27_SIG,
    ROM28_DATA  => ROM21_DATA28_SIG,
    ROM29_DATA  => ROM21_DATA29_SIG,
    ROM30_DATA  => ROM21_DATA30_SIG,
    ROM31_DATA  => ROM21_DATA31_SIG,
    ADDR0       => ADDR21_0_SIG,
    ADDR1       => ADDR21_1_SIG,
    ADDR2       => ADDR21_2_SIG,
    ADDR3       => ADDR21_3_SIG,
    ADDR4       => ADDR21_4_SIG,
    ADDR5       => ADDR21_5_SIG,
    ADDR6       => ADDR21_6_SIG,
    ADDR7       => ADDR21_7_SIG,
    ADDR8       => ADDR21_8_SIG,
    ADDR9       => ADDR21_9_SIG,
    ADDR10      => ADDR21_10_SIG,
    ADDR11      => ADDR21_11_SIG,
    ADDR12      => ADDR21_12_SIG,
    ADDR13      => ADDR21_13_SIG,
    ADDR14      => ADDR21_14_SIG,
    ADDR15      => ADDR21_15_SIG,
    ADDR16      => ADDR21_16_SIG,
    ADDR17      => ADDR21_17_SIG,
    ADDR18      => ADDR21_18_SIG,
    ADDR19      => ADDR21_19_SIG,
    ADDR20      => ADDR21_20_SIG,
    ADDR21      => ADDR21_21_SIG,
    ADDR22      => ADDR21_22_SIG,
    ADDR23      => ADDR21_23_SIG,
    ADDR24      => ADDR21_24_SIG,
    ADDR25      => ADDR21_25_SIG,
    ADDR26      => ADDR21_26_SIG,
    ADDR27      => ADDR21_27_SIG,
    ADDR28      => ADDR21_28_SIG,
    ADDR29      => ADDR21_29_SIG,
    ADDR30      => ADDR21_30_SIG,
    ADDR31      => ADDR21_31_SIG,
    DOUT        => VM21_OUT_SIG
);

VM22_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM22_DATA0_SIG,
    ROM1_DATA   => ROM22_DATA1_SIG,
    ROM2_DATA   => ROM22_DATA2_SIG,
    ROM3_DATA   => ROM22_DATA3_SIG,
    ROM4_DATA   => ROM22_DATA4_SIG,
    ROM5_DATA   => ROM22_DATA5_SIG,
    ROM6_DATA   => ROM22_DATA6_SIG,
    ROM7_DATA   => ROM22_DATA7_SIG,
    ROM8_DATA   => ROM22_DATA8_SIG,
    ROM9_DATA   => ROM22_DATA9_SIG,
    ROM10_DATA  => ROM22_DATA10_SIG,
    ROM11_DATA  => ROM22_DATA11_SIG,
    ROM12_DATA  => ROM22_DATA12_SIG,
    ROM13_DATA  => ROM22_DATA13_SIG,
    ROM14_DATA  => ROM22_DATA14_SIG,
    ROM15_DATA  => ROM22_DATA15_SIG,
    ROM16_DATA  => ROM22_DATA16_SIG,
    ROM17_DATA  => ROM22_DATA17_SIG,
    ROM18_DATA  => ROM22_DATA18_SIG,
    ROM19_DATA  => ROM22_DATA19_SIG,
    ROM20_DATA  => ROM22_DATA20_SIG,
    ROM21_DATA  => ROM22_DATA21_SIG,
    ROM22_DATA  => ROM22_DATA22_SIG,
    ROM23_DATA  => ROM22_DATA23_SIG,
    ROM24_DATA  => ROM22_DATA24_SIG,
    ROM25_DATA  => ROM22_DATA25_SIG,
    ROM26_DATA  => ROM22_DATA26_SIG,
    ROM27_DATA  => ROM22_DATA27_SIG,
    ROM28_DATA  => ROM22_DATA28_SIG,
    ROM29_DATA  => ROM22_DATA29_SIG,
    ROM30_DATA  => ROM22_DATA30_SIG,
    ROM31_DATA  => ROM22_DATA31_SIG,
    ADDR0       => ADDR22_0_SIG,
    ADDR1       => ADDR22_1_SIG,
    ADDR2       => ADDR22_2_SIG,
    ADDR3       => ADDR22_3_SIG,
    ADDR4       => ADDR22_4_SIG,
    ADDR5       => ADDR22_5_SIG,
    ADDR6       => ADDR22_6_SIG,
    ADDR7       => ADDR22_7_SIG,
    ADDR8       => ADDR22_8_SIG,
    ADDR9       => ADDR22_9_SIG,
    ADDR10      => ADDR22_10_SIG,
    ADDR11      => ADDR22_11_SIG,
    ADDR12      => ADDR22_12_SIG,
    ADDR13      => ADDR22_13_SIG,
    ADDR14      => ADDR22_14_SIG,
    ADDR15      => ADDR22_15_SIG,
    ADDR16      => ADDR22_16_SIG,
    ADDR17      => ADDR22_17_SIG,
    ADDR18      => ADDR22_18_SIG,
    ADDR19      => ADDR22_19_SIG,
    ADDR20      => ADDR22_20_SIG,
    ADDR21      => ADDR22_21_SIG,
    ADDR22      => ADDR22_22_SIG,
    ADDR23      => ADDR22_23_SIG,
    ADDR24      => ADDR22_24_SIG,
    ADDR25      => ADDR22_25_SIG,
    ADDR26      => ADDR22_26_SIG,
    ADDR27      => ADDR22_27_SIG,
    ADDR28      => ADDR22_28_SIG,
    ADDR29      => ADDR22_29_SIG,
    ADDR30      => ADDR22_30_SIG,
    ADDR31      => ADDR22_31_SIG,
    DOUT        => VM22_OUT_SIG
);

VM23_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM23_DATA0_SIG,
    ROM1_DATA   => ROM23_DATA1_SIG,
    ROM2_DATA   => ROM23_DATA2_SIG,
    ROM3_DATA   => ROM23_DATA3_SIG,
    ROM4_DATA   => ROM23_DATA4_SIG,
    ROM5_DATA   => ROM23_DATA5_SIG,
    ROM6_DATA   => ROM23_DATA6_SIG,
    ROM7_DATA   => ROM23_DATA7_SIG,
    ROM8_DATA   => ROM23_DATA8_SIG,
    ROM9_DATA   => ROM23_DATA9_SIG,
    ROM10_DATA  => ROM23_DATA10_SIG,
    ROM11_DATA  => ROM23_DATA11_SIG,
    ROM12_DATA  => ROM23_DATA12_SIG,
    ROM13_DATA  => ROM23_DATA13_SIG,
    ROM14_DATA  => ROM23_DATA14_SIG,
    ROM15_DATA  => ROM23_DATA15_SIG,
    ROM16_DATA  => ROM23_DATA16_SIG,
    ROM17_DATA  => ROM23_DATA17_SIG,
    ROM18_DATA  => ROM23_DATA18_SIG,
    ROM19_DATA  => ROM23_DATA19_SIG,
    ROM20_DATA  => ROM23_DATA20_SIG,
    ROM21_DATA  => ROM23_DATA21_SIG,
    ROM22_DATA  => ROM23_DATA22_SIG,
    ROM23_DATA  => ROM23_DATA23_SIG,
    ROM24_DATA  => ROM23_DATA24_SIG,
    ROM25_DATA  => ROM23_DATA25_SIG,
    ROM26_DATA  => ROM23_DATA26_SIG,
    ROM27_DATA  => ROM23_DATA27_SIG,
    ROM28_DATA  => ROM23_DATA28_SIG,
    ROM29_DATA  => ROM23_DATA29_SIG,
    ROM30_DATA  => ROM23_DATA30_SIG,
    ROM31_DATA  => ROM23_DATA31_SIG,
    ADDR0       => ADDR23_0_SIG,
    ADDR1       => ADDR23_1_SIG,
    ADDR2       => ADDR23_2_SIG,
    ADDR3       => ADDR23_3_SIG,
    ADDR4       => ADDR23_4_SIG,
    ADDR5       => ADDR23_5_SIG,
    ADDR6       => ADDR23_6_SIG,
    ADDR7       => ADDR23_7_SIG,
    ADDR8       => ADDR23_8_SIG,
    ADDR9       => ADDR23_9_SIG,
    ADDR10      => ADDR23_10_SIG,
    ADDR11      => ADDR23_11_SIG,
    ADDR12      => ADDR23_12_SIG,
    ADDR13      => ADDR23_13_SIG,
    ADDR14      => ADDR23_14_SIG,
    ADDR15      => ADDR23_15_SIG,
    ADDR16      => ADDR23_16_SIG,
    ADDR17      => ADDR23_17_SIG,
    ADDR18      => ADDR23_18_SIG,
    ADDR19      => ADDR23_19_SIG,
    ADDR20      => ADDR23_20_SIG,
    ADDR21      => ADDR23_21_SIG,
    ADDR22      => ADDR23_22_SIG,
    ADDR23      => ADDR23_23_SIG,
    ADDR24      => ADDR23_24_SIG,
    ADDR25      => ADDR23_25_SIG,
    ADDR26      => ADDR23_26_SIG,
    ADDR27      => ADDR23_27_SIG,
    ADDR28      => ADDR23_28_SIG,
    ADDR29      => ADDR23_29_SIG,
    ADDR30      => ADDR23_30_SIG,
    ADDR31      => ADDR23_31_SIG,
    DOUT        => VM23_OUT_SIG
);

VM24_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM24_DATA0_SIG,
    ROM1_DATA   => ROM24_DATA1_SIG,
    ROM2_DATA   => ROM24_DATA2_SIG,
    ROM3_DATA   => ROM24_DATA3_SIG,
    ROM4_DATA   => ROM24_DATA4_SIG,
    ROM5_DATA   => ROM24_DATA5_SIG,
    ROM6_DATA   => ROM24_DATA6_SIG,
    ROM7_DATA   => ROM24_DATA7_SIG,
    ROM8_DATA   => ROM24_DATA8_SIG,
    ROM9_DATA   => ROM24_DATA9_SIG,
    ROM10_DATA  => ROM24_DATA10_SIG,
    ROM11_DATA  => ROM24_DATA11_SIG,
    ROM12_DATA  => ROM24_DATA12_SIG,
    ROM13_DATA  => ROM24_DATA13_SIG,
    ROM14_DATA  => ROM24_DATA14_SIG,
    ROM15_DATA  => ROM24_DATA15_SIG,
    ROM16_DATA  => ROM24_DATA16_SIG,
    ROM17_DATA  => ROM24_DATA17_SIG,
    ROM18_DATA  => ROM24_DATA18_SIG,
    ROM19_DATA  => ROM24_DATA19_SIG,
    ROM20_DATA  => ROM24_DATA20_SIG,
    ROM21_DATA  => ROM24_DATA21_SIG,
    ROM22_DATA  => ROM24_DATA22_SIG,
    ROM23_DATA  => ROM24_DATA23_SIG,
    ROM24_DATA  => ROM24_DATA24_SIG,
    ROM25_DATA  => ROM24_DATA25_SIG,
    ROM26_DATA  => ROM24_DATA26_SIG,
    ROM27_DATA  => ROM24_DATA27_SIG,
    ROM28_DATA  => ROM24_DATA28_SIG,
    ROM29_DATA  => ROM24_DATA29_SIG,
    ROM30_DATA  => ROM24_DATA30_SIG,
    ROM31_DATA  => ROM24_DATA31_SIG,
    ADDR0       => ADDR24_0_SIG,
    ADDR1       => ADDR24_1_SIG,
    ADDR2       => ADDR24_2_SIG,
    ADDR3       => ADDR24_3_SIG,
    ADDR4       => ADDR24_4_SIG,
    ADDR5       => ADDR24_5_SIG,
    ADDR6       => ADDR24_6_SIG,
    ADDR7       => ADDR24_7_SIG,
    ADDR8       => ADDR24_8_SIG,
    ADDR9       => ADDR24_9_SIG,
    ADDR10      => ADDR24_10_SIG,
    ADDR11      => ADDR24_11_SIG,
    ADDR12      => ADDR24_12_SIG,
    ADDR13      => ADDR24_13_SIG,
    ADDR14      => ADDR24_14_SIG,
    ADDR15      => ADDR24_15_SIG,
    ADDR16      => ADDR24_16_SIG,
    ADDR17      => ADDR24_17_SIG,
    ADDR18      => ADDR24_18_SIG,
    ADDR19      => ADDR24_19_SIG,
    ADDR20      => ADDR24_20_SIG,
    ADDR21      => ADDR24_21_SIG,
    ADDR22      => ADDR24_22_SIG,
    ADDR23      => ADDR24_23_SIG,
    ADDR24      => ADDR24_24_SIG,
    ADDR25      => ADDR24_25_SIG,
    ADDR26      => ADDR24_26_SIG,
    ADDR27      => ADDR24_27_SIG,
    ADDR28      => ADDR24_28_SIG,
    ADDR29      => ADDR24_29_SIG,
    ADDR30      => ADDR24_30_SIG,
    ADDR31      => ADDR24_31_SIG,
    DOUT        => VM24_OUT_SIG
);

VM25_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM25_DATA0_SIG,
    ROM1_DATA   => ROM25_DATA1_SIG,
    ROM2_DATA   => ROM25_DATA2_SIG,
    ROM3_DATA   => ROM25_DATA3_SIG,
    ROM4_DATA   => ROM25_DATA4_SIG,
    ROM5_DATA   => ROM25_DATA5_SIG,
    ROM6_DATA   => ROM25_DATA6_SIG,
    ROM7_DATA   => ROM25_DATA7_SIG,
    ROM8_DATA   => ROM25_DATA8_SIG,
    ROM9_DATA   => ROM25_DATA9_SIG,
    ROM10_DATA  => ROM25_DATA10_SIG,
    ROM11_DATA  => ROM25_DATA11_SIG,
    ROM12_DATA  => ROM25_DATA12_SIG,
    ROM13_DATA  => ROM25_DATA13_SIG,
    ROM14_DATA  => ROM25_DATA14_SIG,
    ROM15_DATA  => ROM25_DATA15_SIG,
    ROM16_DATA  => ROM25_DATA16_SIG,
    ROM17_DATA  => ROM25_DATA17_SIG,
    ROM18_DATA  => ROM25_DATA18_SIG,
    ROM19_DATA  => ROM25_DATA19_SIG,
    ROM20_DATA  => ROM25_DATA20_SIG,
    ROM21_DATA  => ROM25_DATA21_SIG,
    ROM22_DATA  => ROM25_DATA22_SIG,
    ROM23_DATA  => ROM25_DATA23_SIG,
    ROM24_DATA  => ROM25_DATA24_SIG,
    ROM25_DATA  => ROM25_DATA25_SIG,
    ROM26_DATA  => ROM25_DATA26_SIG,
    ROM27_DATA  => ROM25_DATA27_SIG,
    ROM28_DATA  => ROM25_DATA28_SIG,
    ROM29_DATA  => ROM25_DATA29_SIG,
    ROM30_DATA  => ROM25_DATA30_SIG,
    ROM31_DATA  => ROM25_DATA31_SIG,
    ADDR0       => ADDR25_0_SIG,
    ADDR1       => ADDR25_1_SIG,
    ADDR2       => ADDR25_2_SIG,
    ADDR3       => ADDR25_3_SIG,
    ADDR4       => ADDR25_4_SIG,
    ADDR5       => ADDR25_5_SIG,
    ADDR6       => ADDR25_6_SIG,
    ADDR7       => ADDR25_7_SIG,
    ADDR8       => ADDR25_8_SIG,
    ADDR9       => ADDR25_9_SIG,
    ADDR10      => ADDR25_10_SIG,
    ADDR11      => ADDR25_11_SIG,
    ADDR12      => ADDR25_12_SIG,
    ADDR13      => ADDR25_13_SIG,
    ADDR14      => ADDR25_14_SIG,
    ADDR15      => ADDR25_15_SIG,
    ADDR16      => ADDR25_16_SIG,
    ADDR17      => ADDR25_17_SIG,
    ADDR18      => ADDR25_18_SIG,
    ADDR19      => ADDR25_19_SIG,
    ADDR20      => ADDR25_20_SIG,
    ADDR21      => ADDR25_21_SIG,
    ADDR22      => ADDR25_22_SIG,
    ADDR23      => ADDR25_23_SIG,
    ADDR24      => ADDR25_24_SIG,
    ADDR25      => ADDR25_25_SIG,
    ADDR26      => ADDR25_26_SIG,
    ADDR27      => ADDR25_27_SIG,
    ADDR28      => ADDR25_28_SIG,
    ADDR29      => ADDR25_29_SIG,
    ADDR30      => ADDR25_30_SIG,
    ADDR31      => ADDR25_31_SIG,
    DOUT        => VM25_OUT_SIG
);

VM26_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM26_DATA0_SIG,
    ROM1_DATA   => ROM26_DATA1_SIG,
    ROM2_DATA   => ROM26_DATA2_SIG,
    ROM3_DATA   => ROM26_DATA3_SIG,
    ROM4_DATA   => ROM26_DATA4_SIG,
    ROM5_DATA   => ROM26_DATA5_SIG,
    ROM6_DATA   => ROM26_DATA6_SIG,
    ROM7_DATA   => ROM26_DATA7_SIG,
    ROM8_DATA   => ROM26_DATA8_SIG,
    ROM9_DATA   => ROM26_DATA9_SIG,
    ROM10_DATA  => ROM26_DATA10_SIG,
    ROM11_DATA  => ROM26_DATA11_SIG,
    ROM12_DATA  => ROM26_DATA12_SIG,
    ROM13_DATA  => ROM26_DATA13_SIG,
    ROM14_DATA  => ROM26_DATA14_SIG,
    ROM15_DATA  => ROM26_DATA15_SIG,
    ROM16_DATA  => ROM26_DATA16_SIG,
    ROM17_DATA  => ROM26_DATA17_SIG,
    ROM18_DATA  => ROM26_DATA18_SIG,
    ROM19_DATA  => ROM26_DATA19_SIG,
    ROM20_DATA  => ROM26_DATA20_SIG,
    ROM21_DATA  => ROM26_DATA21_SIG,
    ROM22_DATA  => ROM26_DATA22_SIG,
    ROM23_DATA  => ROM26_DATA23_SIG,
    ROM24_DATA  => ROM26_DATA24_SIG,
    ROM25_DATA  => ROM26_DATA25_SIG,
    ROM26_DATA  => ROM26_DATA26_SIG,
    ROM27_DATA  => ROM26_DATA27_SIG,
    ROM28_DATA  => ROM26_DATA28_SIG,
    ROM29_DATA  => ROM26_DATA29_SIG,
    ROM30_DATA  => ROM26_DATA30_SIG,
    ROM31_DATA  => ROM26_DATA31_SIG,
    ADDR0       => ADDR26_0_SIG,
    ADDR1       => ADDR26_1_SIG,
    ADDR2       => ADDR26_2_SIG,
    ADDR3       => ADDR26_3_SIG,
    ADDR4       => ADDR26_4_SIG,
    ADDR5       => ADDR26_5_SIG,
    ADDR6       => ADDR26_6_SIG,
    ADDR7       => ADDR26_7_SIG,
    ADDR8       => ADDR26_8_SIG,
    ADDR9       => ADDR26_9_SIG,
    ADDR10      => ADDR26_10_SIG,
    ADDR11      => ADDR26_11_SIG,
    ADDR12      => ADDR26_12_SIG,
    ADDR13      => ADDR26_13_SIG,
    ADDR14      => ADDR26_14_SIG,
    ADDR15      => ADDR26_15_SIG,
    ADDR16      => ADDR26_16_SIG,
    ADDR17      => ADDR26_17_SIG,
    ADDR18      => ADDR26_18_SIG,
    ADDR19      => ADDR26_19_SIG,
    ADDR20      => ADDR26_20_SIG,
    ADDR21      => ADDR26_21_SIG,
    ADDR22      => ADDR26_22_SIG,
    ADDR23      => ADDR26_23_SIG,
    ADDR24      => ADDR26_24_SIG,
    ADDR25      => ADDR26_25_SIG,
    ADDR26      => ADDR26_26_SIG,
    ADDR27      => ADDR26_27_SIG,
    ADDR28      => ADDR26_28_SIG,
    ADDR29      => ADDR26_29_SIG,
    ADDR30      => ADDR26_30_SIG,
    ADDR31      => ADDR26_31_SIG,
    DOUT        => VM26_OUT_SIG
);

VM27_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM27_DATA0_SIG,
    ROM1_DATA   => ROM27_DATA1_SIG,
    ROM2_DATA   => ROM27_DATA2_SIG,
    ROM3_DATA   => ROM27_DATA3_SIG,
    ROM4_DATA   => ROM27_DATA4_SIG,
    ROM5_DATA   => ROM27_DATA5_SIG,
    ROM6_DATA   => ROM27_DATA6_SIG,
    ROM7_DATA   => ROM27_DATA7_SIG,
    ROM8_DATA   => ROM27_DATA8_SIG,
    ROM9_DATA   => ROM27_DATA9_SIG,
    ROM10_DATA  => ROM27_DATA10_SIG,
    ROM11_DATA  => ROM27_DATA11_SIG,
    ROM12_DATA  => ROM27_DATA12_SIG,
    ROM13_DATA  => ROM27_DATA13_SIG,
    ROM14_DATA  => ROM27_DATA14_SIG,
    ROM15_DATA  => ROM27_DATA15_SIG,
    ROM16_DATA  => ROM27_DATA16_SIG,
    ROM17_DATA  => ROM27_DATA17_SIG,
    ROM18_DATA  => ROM27_DATA18_SIG,
    ROM19_DATA  => ROM27_DATA19_SIG,
    ROM20_DATA  => ROM27_DATA20_SIG,
    ROM21_DATA  => ROM27_DATA21_SIG,
    ROM22_DATA  => ROM27_DATA22_SIG,
    ROM23_DATA  => ROM27_DATA23_SIG,
    ROM24_DATA  => ROM27_DATA24_SIG,
    ROM25_DATA  => ROM27_DATA25_SIG,
    ROM26_DATA  => ROM27_DATA26_SIG,
    ROM27_DATA  => ROM27_DATA27_SIG,
    ROM28_DATA  => ROM27_DATA28_SIG,
    ROM29_DATA  => ROM27_DATA29_SIG,
    ROM30_DATA  => ROM27_DATA30_SIG,
    ROM31_DATA  => ROM27_DATA31_SIG,
    ADDR0       => ADDR27_0_SIG,
    ADDR1       => ADDR27_1_SIG,
    ADDR2       => ADDR27_2_SIG,
    ADDR3       => ADDR27_3_SIG,
    ADDR4       => ADDR27_4_SIG,
    ADDR5       => ADDR27_5_SIG,
    ADDR6       => ADDR27_6_SIG,
    ADDR7       => ADDR27_7_SIG,
    ADDR8       => ADDR27_8_SIG,
    ADDR9       => ADDR27_9_SIG,
    ADDR10      => ADDR27_10_SIG,
    ADDR11      => ADDR27_11_SIG,
    ADDR12      => ADDR27_12_SIG,
    ADDR13      => ADDR27_13_SIG,
    ADDR14      => ADDR27_14_SIG,
    ADDR15      => ADDR27_15_SIG,
    ADDR16      => ADDR27_16_SIG,
    ADDR17      => ADDR27_17_SIG,
    ADDR18      => ADDR27_18_SIG,
    ADDR19      => ADDR27_19_SIG,
    ADDR20      => ADDR27_20_SIG,
    ADDR21      => ADDR27_21_SIG,
    ADDR22      => ADDR27_22_SIG,
    ADDR23      => ADDR27_23_SIG,
    ADDR24      => ADDR27_24_SIG,
    ADDR25      => ADDR27_25_SIG,
    ADDR26      => ADDR27_26_SIG,
    ADDR27      => ADDR27_27_SIG,
    ADDR28      => ADDR27_28_SIG,
    ADDR29      => ADDR27_29_SIG,
    ADDR30      => ADDR27_30_SIG,
    ADDR31      => ADDR27_31_SIG,
    DOUT        => VM27_OUT_SIG
);

VM28_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM28_DATA0_SIG,
    ROM1_DATA   => ROM28_DATA1_SIG,
    ROM2_DATA   => ROM28_DATA2_SIG,
    ROM3_DATA   => ROM28_DATA3_SIG,
    ROM4_DATA   => ROM28_DATA4_SIG,
    ROM5_DATA   => ROM28_DATA5_SIG,
    ROM6_DATA   => ROM28_DATA6_SIG,
    ROM7_DATA   => ROM28_DATA7_SIG,
    ROM8_DATA   => ROM28_DATA8_SIG,
    ROM9_DATA   => ROM28_DATA9_SIG,
    ROM10_DATA  => ROM28_DATA10_SIG,
    ROM11_DATA  => ROM28_DATA11_SIG,
    ROM12_DATA  => ROM28_DATA12_SIG,
    ROM13_DATA  => ROM28_DATA13_SIG,
    ROM14_DATA  => ROM28_DATA14_SIG,
    ROM15_DATA  => ROM28_DATA15_SIG,
    ROM16_DATA  => ROM28_DATA16_SIG,
    ROM17_DATA  => ROM28_DATA17_SIG,
    ROM18_DATA  => ROM28_DATA18_SIG,
    ROM19_DATA  => ROM28_DATA19_SIG,
    ROM20_DATA  => ROM28_DATA20_SIG,
    ROM21_DATA  => ROM28_DATA21_SIG,
    ROM22_DATA  => ROM28_DATA22_SIG,
    ROM23_DATA  => ROM28_DATA23_SIG,
    ROM24_DATA  => ROM28_DATA24_SIG,
    ROM25_DATA  => ROM28_DATA25_SIG,
    ROM26_DATA  => ROM28_DATA26_SIG,
    ROM27_DATA  => ROM28_DATA27_SIG,
    ROM28_DATA  => ROM28_DATA28_SIG,
    ROM29_DATA  => ROM28_DATA29_SIG,
    ROM30_DATA  => ROM28_DATA30_SIG,
    ROM31_DATA  => ROM28_DATA31_SIG,
    ADDR0       => ADDR28_0_SIG,
    ADDR1       => ADDR28_1_SIG,
    ADDR2       => ADDR28_2_SIG,
    ADDR3       => ADDR28_3_SIG,
    ADDR4       => ADDR28_4_SIG,
    ADDR5       => ADDR28_5_SIG,
    ADDR6       => ADDR28_6_SIG,
    ADDR7       => ADDR28_7_SIG,
    ADDR8       => ADDR28_8_SIG,
    ADDR9       => ADDR28_9_SIG,
    ADDR10      => ADDR28_10_SIG,
    ADDR11      => ADDR28_11_SIG,
    ADDR12      => ADDR28_12_SIG,
    ADDR13      => ADDR28_13_SIG,
    ADDR14      => ADDR28_14_SIG,
    ADDR15      => ADDR28_15_SIG,
    ADDR16      => ADDR28_16_SIG,
    ADDR17      => ADDR28_17_SIG,
    ADDR18      => ADDR28_18_SIG,
    ADDR19      => ADDR28_19_SIG,
    ADDR20      => ADDR28_20_SIG,
    ADDR21      => ADDR28_21_SIG,
    ADDR22      => ADDR28_22_SIG,
    ADDR23      => ADDR28_23_SIG,
    ADDR24      => ADDR28_24_SIG,
    ADDR25      => ADDR28_25_SIG,
    ADDR26      => ADDR28_26_SIG,
    ADDR27      => ADDR28_27_SIG,
    ADDR28      => ADDR28_28_SIG,
    ADDR29      => ADDR28_29_SIG,
    ADDR30      => ADDR28_30_SIG,
    ADDR31      => ADDR28_31_SIG,
    DOUT        => VM28_OUT_SIG
);

VM29_INST: VECTOR_MULTIPLIER
Generic map ( WIDTH => 32, POWER =>13 )
Port map (
    CLK         => CLK,
    RESET       => RESET,
    SET         => SET_VM_SIG,
    DIN0        => DIN0_SIG,
    DIN1        => DIN1_SIG,
    DIN2        => DIN2_SIG,
    DIN3        => DIN3_SIG,
    DIN4        => DIN4_SIG,
    DIN5        => DIN5_SIG,
    DIN6        => DIN6_SIG,
    DIN7        => DIN7_SIG,
    DIN8        => DIN8_SIG,
    DIN9        => DIN9_SIG,
    DIN10       => DIN10_SIG,
    DIN11       => DIN11_SIG,
    DIN12       => DIN12_SIG,
    DIN13       => DIN13_SIG,
    DIN14       => DIN14_SIG,
    DIN15       => DIN15_SIG,
    DIN16       => DIN16_SIG,
    DIN17       => DIN17_SIG,
    DIN18       => DIN18_SIG,
    DIN19       => DIN19_SIG,
    DIN20       => DIN20_SIG,
    DIN21       => DIN21_SIG,
    DIN22       => DIN22_SIG,
    DIN23       => DIN23_SIG,
    DIN24       => DIN24_SIG,
    DIN25       => DIN25_SIG,
    DIN26       => DIN26_SIG,
    DIN27       => DIN27_SIG,
    DIN28       => DIN28_SIG,
    DIN29       => DIN29_SIG,
    DIN30       => DIN30_SIG,
    DIN31       => DIN31_SIG,
    ROM0_DATA   => ROM29_DATA0_SIG,
    ROM1_DATA   => ROM29_DATA1_SIG,
    ROM2_DATA   => ROM29_DATA2_SIG,
    ROM3_DATA   => ROM29_DATA3_SIG,
    ROM4_DATA   => ROM29_DATA4_SIG,
    ROM5_DATA   => ROM29_DATA5_SIG,
    ROM6_DATA   => ROM29_DATA6_SIG,
    ROM7_DATA   => ROM29_DATA7_SIG,
    ROM8_DATA   => ROM29_DATA8_SIG,
    ROM9_DATA   => ROM29_DATA9_SIG,
    ROM10_DATA  => ROM29_DATA10_SIG,
    ROM11_DATA  => ROM29_DATA11_SIG,
    ROM12_DATA  => ROM29_DATA12_SIG,
    ROM13_DATA  => ROM29_DATA13_SIG,
    ROM14_DATA  => ROM29_DATA14_SIG,
    ROM15_DATA  => ROM29_DATA15_SIG,
    ROM16_DATA  => ROM29_DATA16_SIG,
    ROM17_DATA  => ROM29_DATA17_SIG,
    ROM18_DATA  => ROM29_DATA18_SIG,
    ROM19_DATA  => ROM29_DATA19_SIG,
    ROM20_DATA  => ROM29_DATA20_SIG,
    ROM21_DATA  => ROM29_DATA21_SIG,
    ROM22_DATA  => ROM29_DATA22_SIG,
    ROM23_DATA  => ROM29_DATA23_SIG,
    ROM24_DATA  => ROM29_DATA24_SIG,
    ROM25_DATA  => ROM29_DATA25_SIG,
    ROM26_DATA  => ROM29_DATA26_SIG,
    ROM27_DATA  => ROM29_DATA27_SIG,
    ROM28_DATA  => ROM29_DATA28_SIG,
    ROM29_DATA  => ROM29_DATA29_SIG,
    ROM30_DATA  => ROM29_DATA30_SIG,
    ROM31_DATA  => ROM29_DATA31_SIG,
    ADDR0       => ADDR29_0_SIG,
    ADDR1       => ADDR29_1_SIG,
    ADDR2       => ADDR29_2_SIG,
    ADDR3       => ADDR29_3_SIG,
    ADDR4       => ADDR29_4_SIG,
    ADDR5       => ADDR29_5_SIG,
    ADDR6       => ADDR29_6_SIG,
    ADDR7       => ADDR29_7_SIG,
    ADDR8       => ADDR29_8_SIG,
    ADDR9       => ADDR29_9_SIG,
    ADDR10      => ADDR29_10_SIG,
    ADDR11      => ADDR29_11_SIG,
    ADDR12      => ADDR29_12_SIG,
    ADDR13      => ADDR29_13_SIG,
    ADDR14      => ADDR29_14_SIG,
    ADDR15      => ADDR29_15_SIG,
    ADDR16      => ADDR29_16_SIG,
    ADDR17      => ADDR29_17_SIG,
    ADDR18      => ADDR29_18_SIG,
    ADDR19      => ADDR29_19_SIG,
    ADDR20      => ADDR29_20_SIG,
    ADDR21      => ADDR29_21_SIG,
    ADDR22      => ADDR29_22_SIG,
    ADDR23      => ADDR29_23_SIG,
    ADDR24      => ADDR29_24_SIG,
    ADDR25      => ADDR29_25_SIG,
    ADDR26      => ADDR29_26_SIG,
    ADDR27      => ADDR29_27_SIG,
    ADDR28      => ADDR29_28_SIG,
    ADDR29      => ADDR29_29_SIG,
    ADDR30      => ADDR29_30_SIG,
    ADDR31      => ADDR29_31_SIG,
    DOUT        => VM29_OUT_SIG
);

COUNTER_FOR_FC_INST: COUNTER_FOR_FC
Port map (
    CLK   => CLK,
    RESET => RESET,
    SET   => SET_CNT_SIG,
    COUT1 => SET_VM_SIG,
    COUT2 => SET_CNT_OL
);

WEIGHT_ROM0_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR0_0_SIG, 
    ADDR1  => ADDR0_1_SIG,
    ADDR2  => ADDR0_2_SIG,
    ADDR3  => ADDR0_3_SIG,
    ADDR4  => ADDR0_4_SIG,
    ADDR5  => ADDR0_5_SIG,
    ADDR6  => ADDR0_6_SIG,
    ADDR7  => ADDR0_7_SIG,
    ADDR8  => ADDR0_8_SIG,
    ADDR9  => ADDR0_9_SIG,
    ADDR10 => ADDR0_10_SIG,
    ADDR11 => ADDR0_11_SIG,
    ADDR12 => ADDR0_12_SIG,
    ADDR13 => ADDR0_13_SIG,
    ADDR14 => ADDR0_14_SIG,
    ADDR15 => ADDR0_15_SIG,
    ADDR16 => ADDR0_16_SIG,
    ADDR17 => ADDR0_17_SIG,
    ADDR18 => ADDR0_18_SIG,
    ADDR19 => ADDR0_19_SIG,
    ADDR20 => ADDR0_20_SIG,
    ADDR21 => ADDR0_21_SIG,
    ADDR22 => ADDR0_22_SIG,
    ADDR23 => ADDR0_23_SIG,
    ADDR24 => ADDR0_24_SIG,
    ADDR25 => ADDR0_25_SIG,
    ADDR26 => ADDR0_26_SIG,
    ADDR27 => ADDR0_27_SIG,
    ADDR28 => ADDR0_28_SIG,
    ADDR29 => ADDR0_29_SIG,
    ADDR30 => ADDR0_30_SIG,
    ADDR31 => ADDR0_31_SIG,
    DATA0  => ROM0_DATA0_SIG,
    DATA1  => ROM0_DATA1_SIG,
    DATA2  => ROM0_DATA2_SIG,
    DATA3  => ROM0_DATA3_SIG,
    DATA4  => ROM0_DATA4_SIG,
    DATA5  => ROM0_DATA5_SIG,
    DATA6  => ROM0_DATA6_SIG,
    DATA7  => ROM0_DATA7_SIG,
    DATA8  => ROM0_DATA8_SIG,
    DATA9  => ROM0_DATA9_SIG,
    DATA10 => ROM0_DATA10_SIG,
    DATA11 => ROM0_DATA11_SIG,
    DATA12 => ROM0_DATA12_SIG,
    DATA13 => ROM0_DATA13_SIG,
    DATA14 => ROM0_DATA14_SIG,
    DATA15 => ROM0_DATA15_SIG,
    DATA16 => ROM0_DATA16_SIG,
    DATA17 => ROM0_DATA17_SIG,
    DATA18 => ROM0_DATA18_SIG,
    DATA19 => ROM0_DATA19_SIG,
    DATA20 => ROM0_DATA20_SIG,
    DATA21 => ROM0_DATA21_SIG,
    DATA22 => ROM0_DATA22_SIG,
    DATA23 => ROM0_DATA23_SIG,
    DATA24 => ROM0_DATA24_SIG,
    DATA25 => ROM0_DATA25_SIG,
    DATA26 => ROM0_DATA26_SIG,
    DATA27 => ROM0_DATA27_SIG,
    DATA28 => ROM0_DATA28_SIG,
    DATA29 => ROM0_DATA29_SIG,
    DATA30 => ROM0_DATA30_SIG,
    DATA31 => ROM0_DATA31_SIG
);

WEIGHT_ROM1_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR1_0_SIG, 
    ADDR1  => ADDR1_1_SIG,
    ADDR2  => ADDR1_2_SIG,
    ADDR3  => ADDR1_3_SIG,
    ADDR4  => ADDR1_4_SIG,
    ADDR5  => ADDR1_5_SIG,
    ADDR6  => ADDR1_6_SIG,
    ADDR7  => ADDR1_7_SIG,
    ADDR8  => ADDR1_8_SIG,
    ADDR9  => ADDR1_9_SIG,
    ADDR10 => ADDR1_10_SIG,
    ADDR11 => ADDR1_11_SIG,
    ADDR12 => ADDR1_12_SIG,
    ADDR13 => ADDR1_13_SIG,
    ADDR14 => ADDR1_14_SIG,
    ADDR15 => ADDR1_15_SIG,
    ADDR16 => ADDR1_16_SIG,
    ADDR17 => ADDR1_17_SIG,
    ADDR18 => ADDR1_18_SIG,
    ADDR19 => ADDR1_19_SIG,
    ADDR20 => ADDR1_20_SIG,
    ADDR21 => ADDR1_21_SIG,
    ADDR22 => ADDR1_22_SIG,
    ADDR23 => ADDR1_23_SIG,
    ADDR24 => ADDR1_24_SIG,
    ADDR25 => ADDR1_25_SIG,
    ADDR26 => ADDR1_26_SIG,
    ADDR27 => ADDR1_27_SIG,
    ADDR28 => ADDR1_28_SIG,
    ADDR29 => ADDR1_29_SIG,
    ADDR30 => ADDR1_30_SIG,
    ADDR31 => ADDR1_31_SIG,
    DATA0  => ROM1_DATA0_SIG,
    DATA1  => ROM1_DATA1_SIG,
    DATA2  => ROM1_DATA2_SIG,
    DATA3  => ROM1_DATA3_SIG,
    DATA4  => ROM1_DATA4_SIG,
    DATA5  => ROM1_DATA5_SIG,
    DATA6  => ROM1_DATA6_SIG,
    DATA7  => ROM1_DATA7_SIG,
    DATA8  => ROM1_DATA8_SIG,
    DATA9  => ROM1_DATA9_SIG,
    DATA10 => ROM1_DATA10_SIG,
    DATA11 => ROM1_DATA11_SIG,
    DATA12 => ROM1_DATA12_SIG,
    DATA13 => ROM1_DATA13_SIG,
    DATA14 => ROM1_DATA14_SIG,
    DATA15 => ROM1_DATA15_SIG,
    DATA16 => ROM1_DATA16_SIG,
    DATA17 => ROM1_DATA17_SIG,
    DATA18 => ROM1_DATA18_SIG,
    DATA19 => ROM1_DATA19_SIG,
    DATA20 => ROM1_DATA20_SIG,
    DATA21 => ROM1_DATA21_SIG,
    DATA22 => ROM1_DATA22_SIG,
    DATA23 => ROM1_DATA23_SIG,
    DATA24 => ROM1_DATA24_SIG,
    DATA25 => ROM1_DATA25_SIG,
    DATA26 => ROM1_DATA26_SIG,
    DATA27 => ROM1_DATA27_SIG,
    DATA28 => ROM1_DATA28_SIG,
    DATA29 => ROM1_DATA29_SIG,
    DATA30 => ROM1_DATA30_SIG,
    DATA31 => ROM1_DATA31_SIG
);

WEIGHT_ROM2_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR2_0_SIG, 
    ADDR1  => ADDR2_1_SIG,
    ADDR2  => ADDR2_2_SIG,
    ADDR3  => ADDR2_3_SIG,
    ADDR4  => ADDR2_4_SIG,
    ADDR5  => ADDR2_5_SIG,
    ADDR6  => ADDR2_6_SIG,
    ADDR7  => ADDR2_7_SIG,
    ADDR8  => ADDR2_8_SIG,
    ADDR9  => ADDR2_9_SIG,
    ADDR10 => ADDR2_10_SIG,
    ADDR11 => ADDR2_11_SIG,
    ADDR12 => ADDR2_12_SIG,
    ADDR13 => ADDR2_13_SIG,
    ADDR14 => ADDR2_14_SIG,
    ADDR15 => ADDR2_15_SIG,
    ADDR16 => ADDR2_16_SIG,
    ADDR17 => ADDR2_17_SIG,
    ADDR18 => ADDR2_18_SIG,
    ADDR19 => ADDR2_19_SIG,
    ADDR20 => ADDR2_20_SIG,
    ADDR21 => ADDR2_21_SIG,
    ADDR22 => ADDR2_22_SIG,
    ADDR23 => ADDR2_23_SIG,
    ADDR24 => ADDR2_24_SIG,
    ADDR25 => ADDR2_25_SIG,
    ADDR26 => ADDR2_26_SIG,
    ADDR27 => ADDR2_27_SIG,
    ADDR28 => ADDR2_28_SIG,
    ADDR29 => ADDR2_29_SIG,
    ADDR30 => ADDR2_30_SIG,
    ADDR31 => ADDR2_31_SIG,
    DATA0  => ROM2_DATA0_SIG,
    DATA1  => ROM2_DATA1_SIG,
    DATA2  => ROM2_DATA2_SIG,
    DATA3  => ROM2_DATA3_SIG,
    DATA4  => ROM2_DATA4_SIG,
    DATA5  => ROM2_DATA5_SIG,
    DATA6  => ROM2_DATA6_SIG,
    DATA7  => ROM2_DATA7_SIG,
    DATA8  => ROM2_DATA8_SIG,
    DATA9  => ROM2_DATA9_SIG,
    DATA10 => ROM2_DATA10_SIG,
    DATA11 => ROM2_DATA11_SIG,
    DATA12 => ROM2_DATA12_SIG,
    DATA13 => ROM2_DATA13_SIG,
    DATA14 => ROM2_DATA14_SIG,
    DATA15 => ROM2_DATA15_SIG,
    DATA16 => ROM2_DATA16_SIG,
    DATA17 => ROM2_DATA17_SIG,
    DATA18 => ROM2_DATA18_SIG,
    DATA19 => ROM2_DATA19_SIG,
    DATA20 => ROM2_DATA20_SIG,
    DATA21 => ROM2_DATA21_SIG,
    DATA22 => ROM2_DATA22_SIG,
    DATA23 => ROM2_DATA23_SIG,
    DATA24 => ROM2_DATA24_SIG,
    DATA25 => ROM2_DATA25_SIG,
    DATA26 => ROM2_DATA26_SIG,
    DATA27 => ROM2_DATA27_SIG,
    DATA28 => ROM2_DATA28_SIG,
    DATA29 => ROM2_DATA29_SIG,
    DATA30 => ROM2_DATA30_SIG,
    DATA31 => ROM2_DATA31_SIG
);

WEIGHT_ROM3_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR3_0_SIG, 
    ADDR1  => ADDR3_1_SIG,
    ADDR2  => ADDR3_2_SIG,
    ADDR3  => ADDR3_3_SIG,
    ADDR4  => ADDR3_4_SIG,
    ADDR5  => ADDR3_5_SIG,
    ADDR6  => ADDR3_6_SIG,
    ADDR7  => ADDR3_7_SIG,
    ADDR8  => ADDR3_8_SIG,
    ADDR9  => ADDR3_9_SIG,
    ADDR10 => ADDR3_10_SIG,
    ADDR11 => ADDR3_11_SIG,
    ADDR12 => ADDR3_12_SIG,
    ADDR13 => ADDR3_13_SIG,
    ADDR14 => ADDR3_14_SIG,
    ADDR15 => ADDR3_15_SIG,
    ADDR16 => ADDR3_16_SIG,
    ADDR17 => ADDR3_17_SIG,
    ADDR18 => ADDR3_18_SIG,
    ADDR19 => ADDR3_19_SIG,
    ADDR20 => ADDR3_20_SIG,
    ADDR21 => ADDR3_21_SIG,
    ADDR22 => ADDR3_22_SIG,
    ADDR23 => ADDR3_23_SIG,
    ADDR24 => ADDR3_24_SIG,
    ADDR25 => ADDR3_25_SIG,
    ADDR26 => ADDR3_26_SIG,
    ADDR27 => ADDR3_27_SIG,
    ADDR28 => ADDR3_28_SIG,
    ADDR29 => ADDR3_29_SIG,
    ADDR30 => ADDR3_30_SIG,
    ADDR31 => ADDR3_31_SIG,
    DATA0  => ROM3_DATA0_SIG,
    DATA1  => ROM3_DATA1_SIG,
    DATA2  => ROM3_DATA2_SIG,
    DATA3  => ROM3_DATA3_SIG,
    DATA4  => ROM3_DATA4_SIG,
    DATA5  => ROM3_DATA5_SIG,
    DATA6  => ROM3_DATA6_SIG,
    DATA7  => ROM3_DATA7_SIG,
    DATA8  => ROM3_DATA8_SIG,
    DATA9  => ROM3_DATA9_SIG,
    DATA10 => ROM3_DATA10_SIG,
    DATA11 => ROM3_DATA11_SIG,
    DATA12 => ROM3_DATA12_SIG,
    DATA13 => ROM3_DATA13_SIG,
    DATA14 => ROM3_DATA14_SIG,
    DATA15 => ROM3_DATA15_SIG,
    DATA16 => ROM3_DATA16_SIG,
    DATA17 => ROM3_DATA17_SIG,
    DATA18 => ROM3_DATA18_SIG,
    DATA19 => ROM3_DATA19_SIG,
    DATA20 => ROM3_DATA20_SIG,
    DATA21 => ROM3_DATA21_SIG,
    DATA22 => ROM3_DATA22_SIG,
    DATA23 => ROM3_DATA23_SIG,
    DATA24 => ROM3_DATA24_SIG,
    DATA25 => ROM3_DATA25_SIG,
    DATA26 => ROM3_DATA26_SIG,
    DATA27 => ROM3_DATA27_SIG,
    DATA28 => ROM3_DATA28_SIG,
    DATA29 => ROM3_DATA29_SIG,
    DATA30 => ROM3_DATA30_SIG,
    DATA31 => ROM3_DATA31_SIG
);

WEIGHT_ROM4_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR4_0_SIG, 
    ADDR1  => ADDR4_1_SIG,
    ADDR2  => ADDR4_2_SIG,
    ADDR3  => ADDR4_3_SIG,
    ADDR4  => ADDR4_4_SIG,
    ADDR5  => ADDR4_5_SIG,
    ADDR6  => ADDR4_6_SIG,
    ADDR7  => ADDR4_7_SIG,
    ADDR8  => ADDR4_8_SIG,
    ADDR9  => ADDR4_9_SIG,
    ADDR10 => ADDR4_10_SIG,
    ADDR11 => ADDR4_11_SIG,
    ADDR12 => ADDR4_12_SIG,
    ADDR13 => ADDR4_13_SIG,
    ADDR14 => ADDR4_14_SIG,
    ADDR15 => ADDR4_15_SIG,
    ADDR16 => ADDR4_16_SIG,
    ADDR17 => ADDR4_17_SIG,
    ADDR18 => ADDR4_18_SIG,
    ADDR19 => ADDR4_19_SIG,
    ADDR20 => ADDR4_20_SIG,
    ADDR21 => ADDR4_21_SIG,
    ADDR22 => ADDR4_22_SIG,
    ADDR23 => ADDR4_23_SIG,
    ADDR24 => ADDR4_24_SIG,
    ADDR25 => ADDR4_25_SIG,
    ADDR26 => ADDR4_26_SIG,
    ADDR27 => ADDR4_27_SIG,
    ADDR28 => ADDR4_28_SIG,
    ADDR29 => ADDR4_29_SIG,
    ADDR30 => ADDR4_30_SIG,
    ADDR31 => ADDR4_31_SIG,
    DATA0  => ROM4_DATA0_SIG,
    DATA1  => ROM4_DATA1_SIG,
    DATA2  => ROM4_DATA2_SIG,
    DATA3  => ROM4_DATA3_SIG,
    DATA4  => ROM4_DATA4_SIG,
    DATA5  => ROM4_DATA5_SIG,
    DATA6  => ROM4_DATA6_SIG,
    DATA7  => ROM4_DATA7_SIG,
    DATA8  => ROM4_DATA8_SIG,
    DATA9  => ROM4_DATA9_SIG,
    DATA10 => ROM4_DATA10_SIG,
    DATA11 => ROM4_DATA11_SIG,
    DATA12 => ROM4_DATA12_SIG,
    DATA13 => ROM4_DATA13_SIG,
    DATA14 => ROM4_DATA14_SIG,
    DATA15 => ROM4_DATA15_SIG,
    DATA16 => ROM4_DATA16_SIG,
    DATA17 => ROM4_DATA17_SIG,
    DATA18 => ROM4_DATA18_SIG,
    DATA19 => ROM4_DATA19_SIG,
    DATA20 => ROM4_DATA20_SIG,
    DATA21 => ROM4_DATA21_SIG,
    DATA22 => ROM4_DATA22_SIG,
    DATA23 => ROM4_DATA23_SIG,
    DATA24 => ROM4_DATA24_SIG,
    DATA25 => ROM4_DATA25_SIG,
    DATA26 => ROM4_DATA26_SIG,
    DATA27 => ROM4_DATA27_SIG,
    DATA28 => ROM4_DATA28_SIG,
    DATA29 => ROM4_DATA29_SIG,
    DATA30 => ROM4_DATA30_SIG,
    DATA31 => ROM4_DATA31_SIG
);

WEIGHT_ROM5_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR5_0_SIG, 
    ADDR1  => ADDR5_1_SIG,
    ADDR2  => ADDR5_2_SIG,
    ADDR3  => ADDR5_3_SIG,
    ADDR4  => ADDR5_4_SIG,
    ADDR5  => ADDR5_5_SIG,
    ADDR6  => ADDR5_6_SIG,
    ADDR7  => ADDR5_7_SIG,
    ADDR8  => ADDR5_8_SIG,
    ADDR9  => ADDR5_9_SIG,
    ADDR10 => ADDR5_10_SIG,
    ADDR11 => ADDR5_11_SIG,
    ADDR12 => ADDR5_12_SIG,
    ADDR13 => ADDR5_13_SIG,
    ADDR14 => ADDR5_14_SIG,
    ADDR15 => ADDR5_15_SIG,
    ADDR16 => ADDR5_16_SIG,
    ADDR17 => ADDR5_17_SIG,
    ADDR18 => ADDR5_18_SIG,
    ADDR19 => ADDR5_19_SIG,
    ADDR20 => ADDR5_20_SIG,
    ADDR21 => ADDR5_21_SIG,
    ADDR22 => ADDR5_22_SIG,
    ADDR23 => ADDR5_23_SIG,
    ADDR24 => ADDR5_24_SIG,
    ADDR25 => ADDR5_25_SIG,
    ADDR26 => ADDR5_26_SIG,
    ADDR27 => ADDR5_27_SIG,
    ADDR28 => ADDR5_28_SIG,
    ADDR29 => ADDR5_29_SIG,
    ADDR30 => ADDR5_30_SIG,
    ADDR31 => ADDR5_31_SIG,
    DATA0  => ROM5_DATA0_SIG,
    DATA1  => ROM5_DATA1_SIG,
    DATA2  => ROM5_DATA2_SIG,
    DATA3  => ROM5_DATA3_SIG,
    DATA4  => ROM5_DATA4_SIG,
    DATA5  => ROM5_DATA5_SIG,
    DATA6  => ROM5_DATA6_SIG,
    DATA7  => ROM5_DATA7_SIG,
    DATA8  => ROM5_DATA8_SIG,
    DATA9  => ROM5_DATA9_SIG,
    DATA10 => ROM5_DATA10_SIG,
    DATA11 => ROM5_DATA11_SIG,
    DATA12 => ROM5_DATA12_SIG,
    DATA13 => ROM5_DATA13_SIG,
    DATA14 => ROM5_DATA14_SIG,
    DATA15 => ROM5_DATA15_SIG,
    DATA16 => ROM5_DATA16_SIG,
    DATA17 => ROM5_DATA17_SIG,
    DATA18 => ROM5_DATA18_SIG,
    DATA19 => ROM5_DATA19_SIG,
    DATA20 => ROM5_DATA20_SIG,
    DATA21 => ROM5_DATA21_SIG,
    DATA22 => ROM5_DATA22_SIG,
    DATA23 => ROM5_DATA23_SIG,
    DATA24 => ROM5_DATA24_SIG,
    DATA25 => ROM5_DATA25_SIG,
    DATA26 => ROM5_DATA26_SIG,
    DATA27 => ROM5_DATA27_SIG,
    DATA28 => ROM5_DATA28_SIG,
    DATA29 => ROM5_DATA29_SIG,
    DATA30 => ROM5_DATA30_SIG,
    DATA31 => ROM5_DATA31_SIG
);

WEIGHT_ROM6_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR6_0_SIG, 
    ADDR1  => ADDR6_1_SIG,
    ADDR2  => ADDR6_2_SIG,
    ADDR3  => ADDR6_3_SIG,
    ADDR4  => ADDR6_4_SIG,
    ADDR5  => ADDR6_5_SIG,
    ADDR6  => ADDR6_6_SIG,
    ADDR7  => ADDR6_7_SIG,
    ADDR8  => ADDR6_8_SIG,
    ADDR9  => ADDR6_9_SIG,
    ADDR10 => ADDR6_10_SIG,
    ADDR11 => ADDR6_11_SIG,
    ADDR12 => ADDR6_12_SIG,
    ADDR13 => ADDR6_13_SIG,
    ADDR14 => ADDR6_14_SIG,
    ADDR15 => ADDR6_15_SIG,
    ADDR16 => ADDR6_16_SIG,
    ADDR17 => ADDR6_17_SIG,
    ADDR18 => ADDR6_18_SIG,
    ADDR19 => ADDR6_19_SIG,
    ADDR20 => ADDR6_20_SIG,
    ADDR21 => ADDR6_21_SIG,
    ADDR22 => ADDR6_22_SIG,
    ADDR23 => ADDR6_23_SIG,
    ADDR24 => ADDR6_24_SIG,
    ADDR25 => ADDR6_25_SIG,
    ADDR26 => ADDR6_26_SIG,
    ADDR27 => ADDR6_27_SIG,
    ADDR28 => ADDR6_28_SIG,
    ADDR29 => ADDR6_29_SIG,
    ADDR30 => ADDR6_30_SIG,
    ADDR31 => ADDR6_31_SIG,
    DATA0  => ROM6_DATA0_SIG,
    DATA1  => ROM6_DATA1_SIG,
    DATA2  => ROM6_DATA2_SIG,
    DATA3  => ROM6_DATA3_SIG,
    DATA4  => ROM6_DATA4_SIG,
    DATA5  => ROM6_DATA5_SIG,
    DATA6  => ROM6_DATA6_SIG,
    DATA7  => ROM6_DATA7_SIG,
    DATA8  => ROM6_DATA8_SIG,
    DATA9  => ROM6_DATA9_SIG,
    DATA10 => ROM6_DATA10_SIG,
    DATA11 => ROM6_DATA11_SIG,
    DATA12 => ROM6_DATA12_SIG,
    DATA13 => ROM6_DATA13_SIG,
    DATA14 => ROM6_DATA14_SIG,
    DATA15 => ROM6_DATA15_SIG,
    DATA16 => ROM6_DATA16_SIG,
    DATA17 => ROM6_DATA17_SIG,
    DATA18 => ROM6_DATA18_SIG,
    DATA19 => ROM6_DATA19_SIG,
    DATA20 => ROM6_DATA20_SIG,
    DATA21 => ROM6_DATA21_SIG,
    DATA22 => ROM6_DATA22_SIG,
    DATA23 => ROM6_DATA23_SIG,
    DATA24 => ROM6_DATA24_SIG,
    DATA25 => ROM6_DATA25_SIG,
    DATA26 => ROM6_DATA26_SIG,
    DATA27 => ROM6_DATA27_SIG,
    DATA28 => ROM6_DATA28_SIG,
    DATA29 => ROM6_DATA29_SIG,
    DATA30 => ROM6_DATA30_SIG,
    DATA31 => ROM6_DATA31_SIG
);

WEIGHT_ROM7_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR7_0_SIG, 
    ADDR1  => ADDR7_1_SIG,
    ADDR2  => ADDR7_2_SIG,
    ADDR3  => ADDR7_3_SIG,
    ADDR4  => ADDR7_4_SIG,
    ADDR5  => ADDR7_5_SIG,
    ADDR6  => ADDR7_6_SIG,
    ADDR7  => ADDR7_7_SIG,
    ADDR8  => ADDR7_8_SIG,
    ADDR9  => ADDR7_9_SIG,
    ADDR10 => ADDR7_10_SIG,
    ADDR11 => ADDR7_11_SIG,
    ADDR12 => ADDR7_12_SIG,
    ADDR13 => ADDR7_13_SIG,
    ADDR14 => ADDR7_14_SIG,
    ADDR15 => ADDR7_15_SIG,
    ADDR16 => ADDR7_16_SIG,
    ADDR17 => ADDR7_17_SIG,
    ADDR18 => ADDR7_18_SIG,
    ADDR19 => ADDR7_19_SIG,
    ADDR20 => ADDR7_20_SIG,
    ADDR21 => ADDR7_21_SIG,
    ADDR22 => ADDR7_22_SIG,
    ADDR23 => ADDR7_23_SIG,
    ADDR24 => ADDR7_24_SIG,
    ADDR25 => ADDR7_25_SIG,
    ADDR26 => ADDR7_26_SIG,
    ADDR27 => ADDR7_27_SIG,
    ADDR28 => ADDR7_28_SIG,
    ADDR29 => ADDR7_29_SIG,
    ADDR30 => ADDR7_30_SIG,
    ADDR31 => ADDR7_31_SIG,
    DATA0  => ROM7_DATA0_SIG,
    DATA1  => ROM7_DATA1_SIG,
    DATA2  => ROM7_DATA2_SIG,
    DATA3  => ROM7_DATA3_SIG,
    DATA4  => ROM7_DATA4_SIG,
    DATA5  => ROM7_DATA5_SIG,
    DATA6  => ROM7_DATA6_SIG,
    DATA7  => ROM7_DATA7_SIG,
    DATA8  => ROM7_DATA8_SIG,
    DATA9  => ROM7_DATA9_SIG,
    DATA10 => ROM7_DATA10_SIG,
    DATA11 => ROM7_DATA11_SIG,
    DATA12 => ROM7_DATA12_SIG,
    DATA13 => ROM7_DATA13_SIG,
    DATA14 => ROM7_DATA14_SIG,
    DATA15 => ROM7_DATA15_SIG,
    DATA16 => ROM7_DATA16_SIG,
    DATA17 => ROM7_DATA17_SIG,
    DATA18 => ROM7_DATA18_SIG,
    DATA19 => ROM7_DATA19_SIG,
    DATA20 => ROM7_DATA20_SIG,
    DATA21 => ROM7_DATA21_SIG,
    DATA22 => ROM7_DATA22_SIG,
    DATA23 => ROM7_DATA23_SIG,
    DATA24 => ROM7_DATA24_SIG,
    DATA25 => ROM7_DATA25_SIG,
    DATA26 => ROM7_DATA26_SIG,
    DATA27 => ROM7_DATA27_SIG,
    DATA28 => ROM7_DATA28_SIG,
    DATA29 => ROM7_DATA29_SIG,
    DATA30 => ROM7_DATA30_SIG,
    DATA31 => ROM7_DATA31_SIG
);

WEIGHT_ROM8_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR8_0_SIG, 
    ADDR1  => ADDR8_1_SIG,
    ADDR2  => ADDR8_2_SIG,
    ADDR3  => ADDR8_3_SIG,
    ADDR4  => ADDR8_4_SIG,
    ADDR5  => ADDR8_5_SIG,
    ADDR6  => ADDR8_6_SIG,
    ADDR7  => ADDR8_7_SIG,
    ADDR8  => ADDR8_8_SIG,
    ADDR9  => ADDR8_9_SIG,
    ADDR10 => ADDR8_10_SIG,
    ADDR11 => ADDR8_11_SIG,
    ADDR12 => ADDR8_12_SIG,
    ADDR13 => ADDR8_13_SIG,
    ADDR14 => ADDR8_14_SIG,
    ADDR15 => ADDR8_15_SIG,
    ADDR16 => ADDR8_16_SIG,
    ADDR17 => ADDR8_17_SIG,
    ADDR18 => ADDR8_18_SIG,
    ADDR19 => ADDR8_19_SIG,
    ADDR20 => ADDR8_20_SIG,
    ADDR21 => ADDR8_21_SIG,
    ADDR22 => ADDR8_22_SIG,
    ADDR23 => ADDR8_23_SIG,
    ADDR24 => ADDR8_24_SIG,
    ADDR25 => ADDR8_25_SIG,
    ADDR26 => ADDR8_26_SIG,
    ADDR27 => ADDR8_27_SIG,
    ADDR28 => ADDR8_28_SIG,
    ADDR29 => ADDR8_29_SIG,
    ADDR30 => ADDR8_30_SIG,
    ADDR31 => ADDR8_31_SIG,
    DATA0  => ROM8_DATA0_SIG,
    DATA1  => ROM8_DATA1_SIG,
    DATA2  => ROM8_DATA2_SIG,
    DATA3  => ROM8_DATA3_SIG,
    DATA4  => ROM8_DATA4_SIG,
    DATA5  => ROM8_DATA5_SIG,
    DATA6  => ROM8_DATA6_SIG,
    DATA7  => ROM8_DATA7_SIG,
    DATA8  => ROM8_DATA8_SIG,
    DATA9  => ROM8_DATA9_SIG,
    DATA10 => ROM8_DATA10_SIG,
    DATA11 => ROM8_DATA11_SIG,
    DATA12 => ROM8_DATA12_SIG,
    DATA13 => ROM8_DATA13_SIG,
    DATA14 => ROM8_DATA14_SIG,
    DATA15 => ROM8_DATA15_SIG,
    DATA16 => ROM8_DATA16_SIG,
    DATA17 => ROM8_DATA17_SIG,
    DATA18 => ROM8_DATA18_SIG,
    DATA19 => ROM8_DATA19_SIG,
    DATA20 => ROM8_DATA20_SIG,
    DATA21 => ROM8_DATA21_SIG,
    DATA22 => ROM8_DATA22_SIG,
    DATA23 => ROM8_DATA23_SIG,
    DATA24 => ROM8_DATA24_SIG,
    DATA25 => ROM8_DATA25_SIG,
    DATA26 => ROM8_DATA26_SIG,
    DATA27 => ROM8_DATA27_SIG,
    DATA28 => ROM8_DATA28_SIG,
    DATA29 => ROM8_DATA29_SIG,
    DATA30 => ROM8_DATA30_SIG,
    DATA31 => ROM8_DATA31_SIG
);

WEIGHT_ROM9_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR9_0_SIG, 
    ADDR1  => ADDR9_1_SIG,
    ADDR2  => ADDR9_2_SIG,
    ADDR3  => ADDR9_3_SIG,
    ADDR4  => ADDR9_4_SIG,
    ADDR5  => ADDR9_5_SIG,
    ADDR6  => ADDR9_6_SIG,
    ADDR7  => ADDR9_7_SIG,
    ADDR8  => ADDR9_8_SIG,
    ADDR9  => ADDR9_9_SIG,
    ADDR10 => ADDR9_10_SIG,
    ADDR11 => ADDR9_11_SIG,
    ADDR12 => ADDR9_12_SIG,
    ADDR13 => ADDR9_13_SIG,
    ADDR14 => ADDR9_14_SIG,
    ADDR15 => ADDR9_15_SIG,
    ADDR16 => ADDR9_16_SIG,
    ADDR17 => ADDR9_17_SIG,
    ADDR18 => ADDR9_18_SIG,
    ADDR19 => ADDR9_19_SIG,
    ADDR20 => ADDR9_20_SIG,
    ADDR21 => ADDR9_21_SIG,
    ADDR22 => ADDR9_22_SIG,
    ADDR23 => ADDR9_23_SIG,
    ADDR24 => ADDR9_24_SIG,
    ADDR25 => ADDR9_25_SIG,
    ADDR26 => ADDR9_26_SIG,
    ADDR27 => ADDR9_27_SIG,
    ADDR28 => ADDR9_28_SIG,
    ADDR29 => ADDR9_29_SIG,
    ADDR30 => ADDR9_30_SIG,
    ADDR31 => ADDR9_31_SIG,
    DATA0  => ROM9_DATA0_SIG,
    DATA1  => ROM9_DATA1_SIG,
    DATA2  => ROM9_DATA2_SIG,
    DATA3  => ROM9_DATA3_SIG,
    DATA4  => ROM9_DATA4_SIG,
    DATA5  => ROM9_DATA5_SIG,
    DATA6  => ROM9_DATA6_SIG,
    DATA7  => ROM9_DATA7_SIG,
    DATA8  => ROM9_DATA8_SIG,
    DATA9  => ROM9_DATA9_SIG,
    DATA10 => ROM9_DATA10_SIG,
    DATA11 => ROM9_DATA11_SIG,
    DATA12 => ROM9_DATA12_SIG,
    DATA13 => ROM9_DATA13_SIG,
    DATA14 => ROM9_DATA14_SIG,
    DATA15 => ROM9_DATA15_SIG,
    DATA16 => ROM9_DATA16_SIG,
    DATA17 => ROM9_DATA17_SIG,
    DATA18 => ROM9_DATA18_SIG,
    DATA19 => ROM9_DATA19_SIG,
    DATA20 => ROM9_DATA20_SIG,
    DATA21 => ROM9_DATA21_SIG,
    DATA22 => ROM9_DATA22_SIG,
    DATA23 => ROM9_DATA23_SIG,
    DATA24 => ROM9_DATA24_SIG,
    DATA25 => ROM9_DATA25_SIG,
    DATA26 => ROM9_DATA26_SIG,
    DATA27 => ROM9_DATA27_SIG,
    DATA28 => ROM9_DATA28_SIG,
    DATA29 => ROM9_DATA29_SIG,
    DATA30 => ROM9_DATA30_SIG,
    DATA31 => ROM9_DATA31_SIG
);

WEIGHT_ROM10_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR10_0_SIG, 
    ADDR1  => ADDR10_1_SIG,
    ADDR2  => ADDR10_2_SIG,
    ADDR3  => ADDR10_3_SIG,
    ADDR4  => ADDR10_4_SIG,
    ADDR5  => ADDR10_5_SIG,
    ADDR6  => ADDR10_6_SIG,
    ADDR7  => ADDR10_7_SIG,
    ADDR8  => ADDR10_8_SIG,
    ADDR9  => ADDR10_9_SIG,
    ADDR10 => ADDR10_10_SIG,
    ADDR11 => ADDR10_11_SIG,
    ADDR12 => ADDR10_12_SIG,
    ADDR13 => ADDR10_13_SIG,
    ADDR14 => ADDR10_14_SIG,
    ADDR15 => ADDR10_15_SIG,
    ADDR16 => ADDR10_16_SIG,
    ADDR17 => ADDR10_17_SIG,
    ADDR18 => ADDR10_18_SIG,
    ADDR19 => ADDR10_19_SIG,
    ADDR20 => ADDR10_20_SIG,
    ADDR21 => ADDR10_21_SIG,
    ADDR22 => ADDR10_22_SIG,
    ADDR23 => ADDR10_23_SIG,
    ADDR24 => ADDR10_24_SIG,
    ADDR25 => ADDR10_25_SIG,
    ADDR26 => ADDR10_26_SIG,
    ADDR27 => ADDR10_27_SIG,
    ADDR28 => ADDR10_28_SIG,
    ADDR29 => ADDR10_29_SIG,
    ADDR30 => ADDR10_30_SIG,
    ADDR31 => ADDR10_31_SIG,
    DATA0  => ROM10_DATA0_SIG,
    DATA1  => ROM10_DATA1_SIG,
    DATA2  => ROM10_DATA2_SIG,
    DATA3  => ROM10_DATA3_SIG,
    DATA4  => ROM10_DATA4_SIG,
    DATA5  => ROM10_DATA5_SIG,
    DATA6  => ROM10_DATA6_SIG,
    DATA7  => ROM10_DATA7_SIG,
    DATA8  => ROM10_DATA8_SIG,
    DATA9  => ROM10_DATA9_SIG,
    DATA10 => ROM10_DATA10_SIG,
    DATA11 => ROM10_DATA11_SIG,
    DATA12 => ROM10_DATA12_SIG,
    DATA13 => ROM10_DATA13_SIG,
    DATA14 => ROM10_DATA14_SIG,
    DATA15 => ROM10_DATA15_SIG,
    DATA16 => ROM10_DATA16_SIG,
    DATA17 => ROM10_DATA17_SIG,
    DATA18 => ROM10_DATA18_SIG,
    DATA19 => ROM10_DATA19_SIG,
    DATA20 => ROM10_DATA20_SIG,
    DATA21 => ROM10_DATA21_SIG,
    DATA22 => ROM10_DATA22_SIG,
    DATA23 => ROM10_DATA23_SIG,
    DATA24 => ROM10_DATA24_SIG,
    DATA25 => ROM10_DATA25_SIG,
    DATA26 => ROM10_DATA26_SIG,
    DATA27 => ROM10_DATA27_SIG,
    DATA28 => ROM10_DATA28_SIG,
    DATA29 => ROM10_DATA29_SIG,
    DATA30 => ROM10_DATA30_SIG,
    DATA31 => ROM10_DATA31_SIG
);

WEIGHT_ROM11_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR11_0_SIG, 
    ADDR1  => ADDR11_1_SIG,
    ADDR2  => ADDR11_2_SIG,
    ADDR3  => ADDR11_3_SIG,
    ADDR4  => ADDR11_4_SIG,
    ADDR5  => ADDR11_5_SIG,
    ADDR6  => ADDR11_6_SIG,
    ADDR7  => ADDR11_7_SIG,
    ADDR8  => ADDR11_8_SIG,
    ADDR9  => ADDR11_9_SIG,
    ADDR10 => ADDR11_10_SIG,
    ADDR11 => ADDR11_11_SIG,
    ADDR12 => ADDR11_12_SIG,
    ADDR13 => ADDR11_13_SIG,
    ADDR14 => ADDR11_14_SIG,
    ADDR15 => ADDR11_15_SIG,
    ADDR16 => ADDR11_16_SIG,
    ADDR17 => ADDR11_17_SIG,
    ADDR18 => ADDR11_18_SIG,
    ADDR19 => ADDR11_19_SIG,
    ADDR20 => ADDR11_20_SIG,
    ADDR21 => ADDR11_21_SIG,
    ADDR22 => ADDR11_22_SIG,
    ADDR23 => ADDR11_23_SIG,
    ADDR24 => ADDR11_24_SIG,
    ADDR25 => ADDR11_25_SIG,
    ADDR26 => ADDR11_26_SIG,
    ADDR27 => ADDR11_27_SIG,
    ADDR28 => ADDR11_28_SIG,
    ADDR29 => ADDR11_29_SIG,
    ADDR30 => ADDR11_30_SIG,
    ADDR31 => ADDR11_31_SIG,
    DATA0  => ROM11_DATA0_SIG,
    DATA1  => ROM11_DATA1_SIG,
    DATA2  => ROM11_DATA2_SIG,
    DATA3  => ROM11_DATA3_SIG,
    DATA4  => ROM11_DATA4_SIG,
    DATA5  => ROM11_DATA5_SIG,
    DATA6  => ROM11_DATA6_SIG,
    DATA7  => ROM11_DATA7_SIG,
    DATA8  => ROM11_DATA8_SIG,
    DATA9  => ROM11_DATA9_SIG,
    DATA10 => ROM11_DATA10_SIG,
    DATA11 => ROM11_DATA11_SIG,
    DATA12 => ROM11_DATA12_SIG,
    DATA13 => ROM11_DATA13_SIG,
    DATA14 => ROM11_DATA14_SIG,
    DATA15 => ROM11_DATA15_SIG,
    DATA16 => ROM11_DATA16_SIG,
    DATA17 => ROM11_DATA17_SIG,
    DATA18 => ROM11_DATA18_SIG,
    DATA19 => ROM11_DATA19_SIG,
    DATA20 => ROM11_DATA20_SIG,
    DATA21 => ROM11_DATA21_SIG,
    DATA22 => ROM11_DATA22_SIG,
    DATA23 => ROM11_DATA23_SIG,
    DATA24 => ROM11_DATA24_SIG,
    DATA25 => ROM11_DATA25_SIG,
    DATA26 => ROM11_DATA26_SIG,
    DATA27 => ROM11_DATA27_SIG,
    DATA28 => ROM11_DATA28_SIG,
    DATA29 => ROM11_DATA29_SIG,
    DATA30 => ROM11_DATA30_SIG,
    DATA31 => ROM11_DATA31_SIG
);

WEIGHT_ROM12_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR12_0_SIG, 
    ADDR1  => ADDR12_1_SIG,
    ADDR2  => ADDR12_2_SIG,
    ADDR3  => ADDR12_3_SIG,
    ADDR4  => ADDR12_4_SIG,
    ADDR5  => ADDR12_5_SIG,
    ADDR6  => ADDR12_6_SIG,
    ADDR7  => ADDR12_7_SIG,
    ADDR8  => ADDR12_8_SIG,
    ADDR9  => ADDR12_9_SIG,
    ADDR10 => ADDR12_10_SIG,
    ADDR11 => ADDR12_11_SIG,
    ADDR12 => ADDR12_12_SIG,
    ADDR13 => ADDR12_13_SIG,
    ADDR14 => ADDR12_14_SIG,
    ADDR15 => ADDR12_15_SIG,
    ADDR16 => ADDR12_16_SIG,
    ADDR17 => ADDR12_17_SIG,
    ADDR18 => ADDR12_18_SIG,
    ADDR19 => ADDR12_19_SIG,
    ADDR20 => ADDR12_20_SIG,
    ADDR21 => ADDR12_21_SIG,
    ADDR22 => ADDR12_22_SIG,
    ADDR23 => ADDR12_23_SIG,
    ADDR24 => ADDR12_24_SIG,
    ADDR25 => ADDR12_25_SIG,
    ADDR26 => ADDR12_26_SIG,
    ADDR27 => ADDR12_27_SIG,
    ADDR28 => ADDR12_28_SIG,
    ADDR29 => ADDR12_29_SIG,
    ADDR30 => ADDR12_30_SIG,
    ADDR31 => ADDR12_31_SIG,
    DATA0  => ROM12_DATA0_SIG,
    DATA1  => ROM12_DATA1_SIG,
    DATA2  => ROM12_DATA2_SIG,
    DATA3  => ROM12_DATA3_SIG,
    DATA4  => ROM12_DATA4_SIG,
    DATA5  => ROM12_DATA5_SIG,
    DATA6  => ROM12_DATA6_SIG,
    DATA7  => ROM12_DATA7_SIG,
    DATA8  => ROM12_DATA8_SIG,
    DATA9  => ROM12_DATA9_SIG,
    DATA10 => ROM12_DATA10_SIG,
    DATA11 => ROM12_DATA11_SIG,
    DATA12 => ROM12_DATA12_SIG,
    DATA13 => ROM12_DATA13_SIG,
    DATA14 => ROM12_DATA14_SIG,
    DATA15 => ROM12_DATA15_SIG,
    DATA16 => ROM12_DATA16_SIG,
    DATA17 => ROM12_DATA17_SIG,
    DATA18 => ROM12_DATA18_SIG,
    DATA19 => ROM12_DATA19_SIG,
    DATA20 => ROM12_DATA20_SIG,
    DATA21 => ROM12_DATA21_SIG,
    DATA22 => ROM12_DATA22_SIG,
    DATA23 => ROM12_DATA23_SIG,
    DATA24 => ROM12_DATA24_SIG,
    DATA25 => ROM12_DATA25_SIG,
    DATA26 => ROM12_DATA26_SIG,
    DATA27 => ROM12_DATA27_SIG,
    DATA28 => ROM12_DATA28_SIG,
    DATA29 => ROM12_DATA29_SIG,
    DATA30 => ROM12_DATA30_SIG,
    DATA31 => ROM12_DATA31_SIG
);

WEIGHT_ROM13_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR13_0_SIG, 
    ADDR1  => ADDR13_1_SIG,
    ADDR2  => ADDR13_2_SIG,
    ADDR3  => ADDR13_3_SIG,
    ADDR4  => ADDR13_4_SIG,
    ADDR5  => ADDR13_5_SIG,
    ADDR6  => ADDR13_6_SIG,
    ADDR7  => ADDR13_7_SIG,
    ADDR8  => ADDR13_8_SIG,
    ADDR9  => ADDR13_9_SIG,
    ADDR10 => ADDR13_10_SIG,
    ADDR11 => ADDR13_11_SIG,
    ADDR12 => ADDR13_12_SIG,
    ADDR13 => ADDR13_13_SIG,
    ADDR14 => ADDR13_14_SIG,
    ADDR15 => ADDR13_15_SIG,
    ADDR16 => ADDR13_16_SIG,
    ADDR17 => ADDR13_17_SIG,
    ADDR18 => ADDR13_18_SIG,
    ADDR19 => ADDR13_19_SIG,
    ADDR20 => ADDR13_20_SIG,
    ADDR21 => ADDR13_21_SIG,
    ADDR22 => ADDR13_22_SIG,
    ADDR23 => ADDR13_23_SIG,
    ADDR24 => ADDR13_24_SIG,
    ADDR25 => ADDR13_25_SIG,
    ADDR26 => ADDR13_26_SIG,
    ADDR27 => ADDR13_27_SIG,
    ADDR28 => ADDR13_28_SIG,
    ADDR29 => ADDR13_29_SIG,
    ADDR30 => ADDR13_30_SIG,
    ADDR31 => ADDR13_31_SIG,
    DATA0  => ROM13_DATA0_SIG,
    DATA1  => ROM13_DATA1_SIG,
    DATA2  => ROM13_DATA2_SIG,
    DATA3  => ROM13_DATA3_SIG,
    DATA4  => ROM13_DATA4_SIG,
    DATA5  => ROM13_DATA5_SIG,
    DATA6  => ROM13_DATA6_SIG,
    DATA7  => ROM13_DATA7_SIG,
    DATA8  => ROM13_DATA8_SIG,
    DATA9  => ROM13_DATA9_SIG,
    DATA10 => ROM13_DATA10_SIG,
    DATA11 => ROM13_DATA11_SIG,
    DATA12 => ROM13_DATA12_SIG,
    DATA13 => ROM13_DATA13_SIG,
    DATA14 => ROM13_DATA14_SIG,
    DATA15 => ROM13_DATA15_SIG,
    DATA16 => ROM13_DATA16_SIG,
    DATA17 => ROM13_DATA17_SIG,
    DATA18 => ROM13_DATA18_SIG,
    DATA19 => ROM13_DATA19_SIG,
    DATA20 => ROM13_DATA20_SIG,
    DATA21 => ROM13_DATA21_SIG,
    DATA22 => ROM13_DATA22_SIG,
    DATA23 => ROM13_DATA23_SIG,
    DATA24 => ROM13_DATA24_SIG,
    DATA25 => ROM13_DATA25_SIG,
    DATA26 => ROM13_DATA26_SIG,
    DATA27 => ROM13_DATA27_SIG,
    DATA28 => ROM13_DATA28_SIG,
    DATA29 => ROM13_DATA29_SIG,
    DATA30 => ROM13_DATA30_SIG,
    DATA31 => ROM13_DATA31_SIG
);

WEIGHT_ROM14_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR14_0_SIG, 
    ADDR1  => ADDR14_1_SIG,
    ADDR2  => ADDR14_2_SIG,
    ADDR3  => ADDR14_3_SIG,
    ADDR4  => ADDR14_4_SIG,
    ADDR5  => ADDR14_5_SIG,
    ADDR6  => ADDR14_6_SIG,
    ADDR7  => ADDR14_7_SIG,
    ADDR8  => ADDR14_8_SIG,
    ADDR9  => ADDR14_9_SIG,
    ADDR10 => ADDR14_10_SIG,
    ADDR11 => ADDR14_11_SIG,
    ADDR12 => ADDR14_12_SIG,
    ADDR13 => ADDR14_13_SIG,
    ADDR14 => ADDR14_14_SIG,
    ADDR15 => ADDR14_15_SIG,
    ADDR16 => ADDR14_16_SIG,
    ADDR17 => ADDR14_17_SIG,
    ADDR18 => ADDR14_18_SIG,
    ADDR19 => ADDR14_19_SIG,
    ADDR20 => ADDR14_20_SIG,
    ADDR21 => ADDR14_21_SIG,
    ADDR22 => ADDR14_22_SIG,
    ADDR23 => ADDR14_23_SIG,
    ADDR24 => ADDR14_24_SIG,
    ADDR25 => ADDR14_25_SIG,
    ADDR26 => ADDR14_26_SIG,
    ADDR27 => ADDR14_27_SIG,
    ADDR28 => ADDR14_28_SIG,
    ADDR29 => ADDR14_29_SIG,
    ADDR30 => ADDR14_30_SIG,
    ADDR31 => ADDR14_31_SIG,
    DATA0  => ROM14_DATA0_SIG,
    DATA1  => ROM14_DATA1_SIG,
    DATA2  => ROM14_DATA2_SIG,
    DATA3  => ROM14_DATA3_SIG,
    DATA4  => ROM14_DATA4_SIG,
    DATA5  => ROM14_DATA5_SIG,
    DATA6  => ROM14_DATA6_SIG,
    DATA7  => ROM14_DATA7_SIG,
    DATA8  => ROM14_DATA8_SIG,
    DATA9  => ROM14_DATA9_SIG,
    DATA10 => ROM14_DATA10_SIG,
    DATA11 => ROM14_DATA11_SIG,
    DATA12 => ROM14_DATA12_SIG,
    DATA13 => ROM14_DATA13_SIG,
    DATA14 => ROM14_DATA14_SIG,
    DATA15 => ROM14_DATA15_SIG,
    DATA16 => ROM14_DATA16_SIG,
    DATA17 => ROM14_DATA17_SIG,
    DATA18 => ROM14_DATA18_SIG,
    DATA19 => ROM14_DATA19_SIG,
    DATA20 => ROM14_DATA20_SIG,
    DATA21 => ROM14_DATA21_SIG,
    DATA22 => ROM14_DATA22_SIG,
    DATA23 => ROM14_DATA23_SIG,
    DATA24 => ROM14_DATA24_SIG,
    DATA25 => ROM14_DATA25_SIG,
    DATA26 => ROM14_DATA26_SIG,
    DATA27 => ROM14_DATA27_SIG,
    DATA28 => ROM14_DATA28_SIG,
    DATA29 => ROM14_DATA29_SIG,
    DATA30 => ROM14_DATA30_SIG,
    DATA31 => ROM14_DATA31_SIG
);

WEIGHT_ROM15_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR15_0_SIG, 
    ADDR1  => ADDR15_1_SIG,
    ADDR2  => ADDR15_2_SIG,
    ADDR3  => ADDR15_3_SIG,
    ADDR4  => ADDR15_4_SIG,
    ADDR5  => ADDR15_5_SIG,
    ADDR6  => ADDR15_6_SIG,
    ADDR7  => ADDR15_7_SIG,
    ADDR8  => ADDR15_8_SIG,
    ADDR9  => ADDR15_9_SIG,
    ADDR10 => ADDR15_10_SIG,
    ADDR11 => ADDR15_11_SIG,
    ADDR12 => ADDR15_12_SIG,
    ADDR13 => ADDR15_13_SIG,
    ADDR14 => ADDR15_14_SIG,
    ADDR15 => ADDR15_15_SIG,
    ADDR16 => ADDR15_16_SIG,
    ADDR17 => ADDR15_17_SIG,
    ADDR18 => ADDR15_18_SIG,
    ADDR19 => ADDR15_19_SIG,
    ADDR20 => ADDR15_20_SIG,
    ADDR21 => ADDR15_21_SIG,
    ADDR22 => ADDR15_22_SIG,
    ADDR23 => ADDR15_23_SIG,
    ADDR24 => ADDR15_24_SIG,
    ADDR25 => ADDR15_25_SIG,
    ADDR26 => ADDR15_26_SIG,
    ADDR27 => ADDR15_27_SIG,
    ADDR28 => ADDR15_28_SIG,
    ADDR29 => ADDR15_29_SIG,
    ADDR30 => ADDR15_30_SIG,
    ADDR31 => ADDR15_31_SIG,
    DATA0  => ROM15_DATA0_SIG,
    DATA1  => ROM15_DATA1_SIG,
    DATA2  => ROM15_DATA2_SIG,
    DATA3  => ROM15_DATA3_SIG,
    DATA4  => ROM15_DATA4_SIG,
    DATA5  => ROM15_DATA5_SIG,
    DATA6  => ROM15_DATA6_SIG,
    DATA7  => ROM15_DATA7_SIG,
    DATA8  => ROM15_DATA8_SIG,
    DATA9  => ROM15_DATA9_SIG,
    DATA10 => ROM15_DATA10_SIG,
    DATA11 => ROM15_DATA11_SIG,
    DATA12 => ROM15_DATA12_SIG,
    DATA13 => ROM15_DATA13_SIG,
    DATA14 => ROM15_DATA14_SIG,
    DATA15 => ROM15_DATA15_SIG,
    DATA16 => ROM15_DATA16_SIG,
    DATA17 => ROM15_DATA17_SIG,
    DATA18 => ROM15_DATA18_SIG,
    DATA19 => ROM15_DATA19_SIG,
    DATA20 => ROM15_DATA20_SIG,
    DATA21 => ROM15_DATA21_SIG,
    DATA22 => ROM15_DATA22_SIG,
    DATA23 => ROM15_DATA23_SIG,
    DATA24 => ROM15_DATA24_SIG,
    DATA25 => ROM15_DATA25_SIG,
    DATA26 => ROM15_DATA26_SIG,
    DATA27 => ROM15_DATA27_SIG,
    DATA28 => ROM15_DATA28_SIG,
    DATA29 => ROM15_DATA29_SIG,
    DATA30 => ROM15_DATA30_SIG,
    DATA31 => ROM15_DATA31_SIG
);

WEIGHT_ROM16_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR16_0_SIG, 
    ADDR1  => ADDR16_1_SIG,
    ADDR2  => ADDR16_2_SIG,
    ADDR3  => ADDR16_3_SIG,
    ADDR4  => ADDR16_4_SIG,
    ADDR5  => ADDR16_5_SIG,
    ADDR6  => ADDR16_6_SIG,
    ADDR7  => ADDR16_7_SIG,
    ADDR8  => ADDR16_8_SIG,
    ADDR9  => ADDR16_9_SIG,
    ADDR10 => ADDR16_10_SIG,
    ADDR11 => ADDR16_11_SIG,
    ADDR12 => ADDR16_12_SIG,
    ADDR13 => ADDR16_13_SIG,
    ADDR14 => ADDR16_14_SIG,
    ADDR15 => ADDR16_15_SIG,
    ADDR16 => ADDR16_16_SIG,
    ADDR17 => ADDR16_17_SIG,
    ADDR18 => ADDR16_18_SIG,
    ADDR19 => ADDR16_19_SIG,
    ADDR20 => ADDR16_20_SIG,
    ADDR21 => ADDR16_21_SIG,
    ADDR22 => ADDR16_22_SIG,
    ADDR23 => ADDR16_23_SIG,
    ADDR24 => ADDR16_24_SIG,
    ADDR25 => ADDR16_25_SIG,
    ADDR26 => ADDR16_26_SIG,
    ADDR27 => ADDR16_27_SIG,
    ADDR28 => ADDR16_28_SIG,
    ADDR29 => ADDR16_29_SIG,
    ADDR30 => ADDR16_30_SIG,
    ADDR31 => ADDR16_31_SIG,
    DATA0  => ROM16_DATA0_SIG,
    DATA1  => ROM16_DATA1_SIG,
    DATA2  => ROM16_DATA2_SIG,
    DATA3  => ROM16_DATA3_SIG,
    DATA4  => ROM16_DATA4_SIG,
    DATA5  => ROM16_DATA5_SIG,
    DATA6  => ROM16_DATA6_SIG,
    DATA7  => ROM16_DATA7_SIG,
    DATA8  => ROM16_DATA8_SIG,
    DATA9  => ROM16_DATA9_SIG,
    DATA10 => ROM16_DATA10_SIG,
    DATA11 => ROM16_DATA11_SIG,
    DATA12 => ROM16_DATA12_SIG,
    DATA13 => ROM16_DATA13_SIG,
    DATA14 => ROM16_DATA14_SIG,
    DATA15 => ROM16_DATA15_SIG,
    DATA16 => ROM16_DATA16_SIG,
    DATA17 => ROM16_DATA17_SIG,
    DATA18 => ROM16_DATA18_SIG,
    DATA19 => ROM16_DATA19_SIG,
    DATA20 => ROM16_DATA20_SIG,
    DATA21 => ROM16_DATA21_SIG,
    DATA22 => ROM16_DATA22_SIG,
    DATA23 => ROM16_DATA23_SIG,
    DATA24 => ROM16_DATA24_SIG,
    DATA25 => ROM16_DATA25_SIG,
    DATA26 => ROM16_DATA26_SIG,
    DATA27 => ROM16_DATA27_SIG,
    DATA28 => ROM16_DATA28_SIG,
    DATA29 => ROM16_DATA29_SIG,
    DATA30 => ROM16_DATA30_SIG,
    DATA31 => ROM16_DATA31_SIG
);

WEIGHT_ROM17_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR17_0_SIG, 
    ADDR1  => ADDR17_1_SIG,
    ADDR2  => ADDR17_2_SIG,
    ADDR3  => ADDR17_3_SIG,
    ADDR4  => ADDR17_4_SIG,
    ADDR5  => ADDR17_5_SIG,
    ADDR6  => ADDR17_6_SIG,
    ADDR7  => ADDR17_7_SIG,
    ADDR8  => ADDR17_8_SIG,
    ADDR9  => ADDR17_9_SIG,
    ADDR10 => ADDR17_10_SIG,
    ADDR11 => ADDR17_11_SIG,
    ADDR12 => ADDR17_12_SIG,
    ADDR13 => ADDR17_13_SIG,
    ADDR14 => ADDR17_14_SIG,
    ADDR15 => ADDR17_15_SIG,
    ADDR16 => ADDR17_16_SIG,
    ADDR17 => ADDR17_17_SIG,
    ADDR18 => ADDR17_18_SIG,
    ADDR19 => ADDR17_19_SIG,
    ADDR20 => ADDR17_20_SIG,
    ADDR21 => ADDR17_21_SIG,
    ADDR22 => ADDR17_22_SIG,
    ADDR23 => ADDR17_23_SIG,
    ADDR24 => ADDR17_24_SIG,
    ADDR25 => ADDR17_25_SIG,
    ADDR26 => ADDR17_26_SIG,
    ADDR27 => ADDR17_27_SIG,
    ADDR28 => ADDR17_28_SIG,
    ADDR29 => ADDR17_29_SIG,
    ADDR30 => ADDR17_30_SIG,
    ADDR31 => ADDR17_31_SIG,
    DATA0  => ROM17_DATA0_SIG,
    DATA1  => ROM17_DATA1_SIG,
    DATA2  => ROM17_DATA2_SIG,
    DATA3  => ROM17_DATA3_SIG,
    DATA4  => ROM17_DATA4_SIG,
    DATA5  => ROM17_DATA5_SIG,
    DATA6  => ROM17_DATA6_SIG,
    DATA7  => ROM17_DATA7_SIG,
    DATA8  => ROM17_DATA8_SIG,
    DATA9  => ROM17_DATA9_SIG,
    DATA10 => ROM17_DATA10_SIG,
    DATA11 => ROM17_DATA11_SIG,
    DATA12 => ROM17_DATA12_SIG,
    DATA13 => ROM17_DATA13_SIG,
    DATA14 => ROM17_DATA14_SIG,
    DATA15 => ROM17_DATA15_SIG,
    DATA16 => ROM17_DATA16_SIG,
    DATA17 => ROM17_DATA17_SIG,
    DATA18 => ROM17_DATA18_SIG,
    DATA19 => ROM17_DATA19_SIG,
    DATA20 => ROM17_DATA20_SIG,
    DATA21 => ROM17_DATA21_SIG,
    DATA22 => ROM17_DATA22_SIG,
    DATA23 => ROM17_DATA23_SIG,
    DATA24 => ROM17_DATA24_SIG,
    DATA25 => ROM17_DATA25_SIG,
    DATA26 => ROM17_DATA26_SIG,
    DATA27 => ROM17_DATA27_SIG,
    DATA28 => ROM17_DATA28_SIG,
    DATA29 => ROM17_DATA29_SIG,
    DATA30 => ROM17_DATA30_SIG,
    DATA31 => ROM17_DATA31_SIG
);

WEIGHT_ROM18_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR18_0_SIG, 
    ADDR1  => ADDR18_1_SIG,
    ADDR2  => ADDR18_2_SIG,
    ADDR3  => ADDR18_3_SIG,
    ADDR4  => ADDR18_4_SIG,
    ADDR5  => ADDR18_5_SIG,
    ADDR6  => ADDR18_6_SIG,
    ADDR7  => ADDR18_7_SIG,
    ADDR8  => ADDR18_8_SIG,
    ADDR9  => ADDR18_9_SIG,
    ADDR10 => ADDR18_10_SIG,
    ADDR11 => ADDR18_11_SIG,
    ADDR12 => ADDR18_12_SIG,
    ADDR13 => ADDR18_13_SIG,
    ADDR14 => ADDR18_14_SIG,
    ADDR15 => ADDR18_15_SIG,
    ADDR16 => ADDR18_16_SIG,
    ADDR17 => ADDR18_17_SIG,
    ADDR18 => ADDR18_18_SIG,
    ADDR19 => ADDR18_19_SIG,
    ADDR20 => ADDR18_20_SIG,
    ADDR21 => ADDR18_21_SIG,
    ADDR22 => ADDR18_22_SIG,
    ADDR23 => ADDR18_23_SIG,
    ADDR24 => ADDR18_24_SIG,
    ADDR25 => ADDR18_25_SIG,
    ADDR26 => ADDR18_26_SIG,
    ADDR27 => ADDR18_27_SIG,
    ADDR28 => ADDR18_28_SIG,
    ADDR29 => ADDR18_29_SIG,
    ADDR30 => ADDR18_30_SIG,
    ADDR31 => ADDR18_31_SIG,
    DATA0  => ROM18_DATA0_SIG,
    DATA1  => ROM18_DATA1_SIG,
    DATA2  => ROM18_DATA2_SIG,
    DATA3  => ROM18_DATA3_SIG,
    DATA4  => ROM18_DATA4_SIG,
    DATA5  => ROM18_DATA5_SIG,
    DATA6  => ROM18_DATA6_SIG,
    DATA7  => ROM18_DATA7_SIG,
    DATA8  => ROM18_DATA8_SIG,
    DATA9  => ROM18_DATA9_SIG,
    DATA10 => ROM18_DATA10_SIG,
    DATA11 => ROM18_DATA11_SIG,
    DATA12 => ROM18_DATA12_SIG,
    DATA13 => ROM18_DATA13_SIG,
    DATA14 => ROM18_DATA14_SIG,
    DATA15 => ROM18_DATA15_SIG,
    DATA16 => ROM18_DATA16_SIG,
    DATA17 => ROM18_DATA17_SIG,
    DATA18 => ROM18_DATA18_SIG,
    DATA19 => ROM18_DATA19_SIG,
    DATA20 => ROM18_DATA20_SIG,
    DATA21 => ROM18_DATA21_SIG,
    DATA22 => ROM18_DATA22_SIG,
    DATA23 => ROM18_DATA23_SIG,
    DATA24 => ROM18_DATA24_SIG,
    DATA25 => ROM18_DATA25_SIG,
    DATA26 => ROM18_DATA26_SIG,
    DATA27 => ROM18_DATA27_SIG,
    DATA28 => ROM18_DATA28_SIG,
    DATA29 => ROM18_DATA29_SIG,
    DATA30 => ROM18_DATA30_SIG,
    DATA31 => ROM18_DATA31_SIG
);

WEIGHT_ROM19_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR19_0_SIG, 
    ADDR1  => ADDR19_1_SIG,
    ADDR2  => ADDR19_2_SIG,
    ADDR3  => ADDR19_3_SIG,
    ADDR4  => ADDR19_4_SIG,
    ADDR5  => ADDR19_5_SIG,
    ADDR6  => ADDR19_6_SIG,
    ADDR7  => ADDR19_7_SIG,
    ADDR8  => ADDR19_8_SIG,
    ADDR9  => ADDR19_9_SIG,
    ADDR10 => ADDR19_10_SIG,
    ADDR11 => ADDR19_11_SIG,
    ADDR12 => ADDR19_12_SIG,
    ADDR13 => ADDR19_13_SIG,
    ADDR14 => ADDR19_14_SIG,
    ADDR15 => ADDR19_15_SIG,
    ADDR16 => ADDR19_16_SIG,
    ADDR17 => ADDR19_17_SIG,
    ADDR18 => ADDR19_18_SIG,
    ADDR19 => ADDR19_19_SIG,
    ADDR20 => ADDR19_20_SIG,
    ADDR21 => ADDR19_21_SIG,
    ADDR22 => ADDR19_22_SIG,
    ADDR23 => ADDR19_23_SIG,
    ADDR24 => ADDR19_24_SIG,
    ADDR25 => ADDR19_25_SIG,
    ADDR26 => ADDR19_26_SIG,
    ADDR27 => ADDR19_27_SIG,
    ADDR28 => ADDR19_28_SIG,
    ADDR29 => ADDR19_29_SIG,
    ADDR30 => ADDR19_30_SIG,
    ADDR31 => ADDR19_31_SIG,
    DATA0  => ROM19_DATA0_SIG,
    DATA1  => ROM19_DATA1_SIG,
    DATA2  => ROM19_DATA2_SIG,
    DATA3  => ROM19_DATA3_SIG,
    DATA4  => ROM19_DATA4_SIG,
    DATA5  => ROM19_DATA5_SIG,
    DATA6  => ROM19_DATA6_SIG,
    DATA7  => ROM19_DATA7_SIG,
    DATA8  => ROM19_DATA8_SIG,
    DATA9  => ROM19_DATA9_SIG,
    DATA10 => ROM19_DATA10_SIG,
    DATA11 => ROM19_DATA11_SIG,
    DATA12 => ROM19_DATA12_SIG,
    DATA13 => ROM19_DATA13_SIG,
    DATA14 => ROM19_DATA14_SIG,
    DATA15 => ROM19_DATA15_SIG,
    DATA16 => ROM19_DATA16_SIG,
    DATA17 => ROM19_DATA17_SIG,
    DATA18 => ROM19_DATA18_SIG,
    DATA19 => ROM19_DATA19_SIG,
    DATA20 => ROM19_DATA20_SIG,
    DATA21 => ROM19_DATA21_SIG,
    DATA22 => ROM19_DATA22_SIG,
    DATA23 => ROM19_DATA23_SIG,
    DATA24 => ROM19_DATA24_SIG,
    DATA25 => ROM19_DATA25_SIG,
    DATA26 => ROM19_DATA26_SIG,
    DATA27 => ROM19_DATA27_SIG,
    DATA28 => ROM19_DATA28_SIG,
    DATA29 => ROM19_DATA29_SIG,
    DATA30 => ROM19_DATA30_SIG,
    DATA31 => ROM19_DATA31_SIG
);

WEIGHT_ROM20_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR20_0_SIG, 
    ADDR1  => ADDR20_1_SIG,
    ADDR2  => ADDR20_2_SIG,
    ADDR3  => ADDR20_3_SIG,
    ADDR4  => ADDR20_4_SIG,
    ADDR5  => ADDR20_5_SIG,
    ADDR6  => ADDR20_6_SIG,
    ADDR7  => ADDR20_7_SIG,
    ADDR8  => ADDR20_8_SIG,
    ADDR9  => ADDR20_9_SIG,
    ADDR10 => ADDR20_10_SIG,
    ADDR11 => ADDR20_11_SIG,
    ADDR12 => ADDR20_12_SIG,
    ADDR13 => ADDR20_13_SIG,
    ADDR14 => ADDR20_14_SIG,
    ADDR15 => ADDR20_15_SIG,
    ADDR16 => ADDR20_16_SIG,
    ADDR17 => ADDR20_17_SIG,
    ADDR18 => ADDR20_18_SIG,
    ADDR19 => ADDR20_19_SIG,
    ADDR20 => ADDR20_20_SIG,
    ADDR21 => ADDR20_21_SIG,
    ADDR22 => ADDR20_22_SIG,
    ADDR23 => ADDR20_23_SIG,
    ADDR24 => ADDR20_24_SIG,
    ADDR25 => ADDR20_25_SIG,
    ADDR26 => ADDR20_26_SIG,
    ADDR27 => ADDR20_27_SIG,
    ADDR28 => ADDR20_28_SIG,
    ADDR29 => ADDR20_29_SIG,
    ADDR30 => ADDR20_30_SIG,
    ADDR31 => ADDR20_31_SIG,
    DATA0  => ROM20_DATA0_SIG,
    DATA1  => ROM20_DATA1_SIG,
    DATA2  => ROM20_DATA2_SIG,
    DATA3  => ROM20_DATA3_SIG,
    DATA4  => ROM20_DATA4_SIG,
    DATA5  => ROM20_DATA5_SIG,
    DATA6  => ROM20_DATA6_SIG,
    DATA7  => ROM20_DATA7_SIG,
    DATA8  => ROM20_DATA8_SIG,
    DATA9  => ROM20_DATA9_SIG,
    DATA10 => ROM20_DATA10_SIG,
    DATA11 => ROM20_DATA11_SIG,
    DATA12 => ROM20_DATA12_SIG,
    DATA13 => ROM20_DATA13_SIG,
    DATA14 => ROM20_DATA14_SIG,
    DATA15 => ROM20_DATA15_SIG,
    DATA16 => ROM20_DATA16_SIG,
    DATA17 => ROM20_DATA17_SIG,
    DATA18 => ROM20_DATA18_SIG,
    DATA19 => ROM20_DATA19_SIG,
    DATA20 => ROM20_DATA20_SIG,
    DATA21 => ROM20_DATA21_SIG,
    DATA22 => ROM20_DATA22_SIG,
    DATA23 => ROM20_DATA23_SIG,
    DATA24 => ROM20_DATA24_SIG,
    DATA25 => ROM20_DATA25_SIG,
    DATA26 => ROM20_DATA26_SIG,
    DATA27 => ROM20_DATA27_SIG,
    DATA28 => ROM20_DATA28_SIG,
    DATA29 => ROM20_DATA29_SIG,
    DATA30 => ROM20_DATA30_SIG,
    DATA31 => ROM20_DATA31_SIG
);

WEIGHT_ROM21_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR21_0_SIG, 
    ADDR1  => ADDR21_1_SIG,
    ADDR2  => ADDR21_2_SIG,
    ADDR3  => ADDR21_3_SIG,
    ADDR4  => ADDR21_4_SIG,
    ADDR5  => ADDR21_5_SIG,
    ADDR6  => ADDR21_6_SIG,
    ADDR7  => ADDR21_7_SIG,
    ADDR8  => ADDR21_8_SIG,
    ADDR9  => ADDR21_9_SIG,
    ADDR10 => ADDR21_10_SIG,
    ADDR11 => ADDR21_11_SIG,
    ADDR12 => ADDR21_12_SIG,
    ADDR13 => ADDR21_13_SIG,
    ADDR14 => ADDR21_14_SIG,
    ADDR15 => ADDR21_15_SIG,
    ADDR16 => ADDR21_16_SIG,
    ADDR17 => ADDR21_17_SIG,
    ADDR18 => ADDR21_18_SIG,
    ADDR19 => ADDR21_19_SIG,
    ADDR20 => ADDR21_20_SIG,
    ADDR21 => ADDR21_21_SIG,
    ADDR22 => ADDR21_22_SIG,
    ADDR23 => ADDR21_23_SIG,
    ADDR24 => ADDR21_24_SIG,
    ADDR25 => ADDR21_25_SIG,
    ADDR26 => ADDR21_26_SIG,
    ADDR27 => ADDR21_27_SIG,
    ADDR28 => ADDR21_28_SIG,
    ADDR29 => ADDR21_29_SIG,
    ADDR30 => ADDR21_30_SIG,
    ADDR31 => ADDR21_31_SIG,
    DATA0  => ROM21_DATA0_SIG,
    DATA1  => ROM21_DATA1_SIG,
    DATA2  => ROM21_DATA2_SIG,
    DATA3  => ROM21_DATA3_SIG,
    DATA4  => ROM21_DATA4_SIG,
    DATA5  => ROM21_DATA5_SIG,
    DATA6  => ROM21_DATA6_SIG,
    DATA7  => ROM21_DATA7_SIG,
    DATA8  => ROM21_DATA8_SIG,
    DATA9  => ROM21_DATA9_SIG,
    DATA10 => ROM21_DATA10_SIG,
    DATA11 => ROM21_DATA11_SIG,
    DATA12 => ROM21_DATA12_SIG,
    DATA13 => ROM21_DATA13_SIG,
    DATA14 => ROM21_DATA14_SIG,
    DATA15 => ROM21_DATA15_SIG,
    DATA16 => ROM21_DATA16_SIG,
    DATA17 => ROM21_DATA17_SIG,
    DATA18 => ROM21_DATA18_SIG,
    DATA19 => ROM21_DATA19_SIG,
    DATA20 => ROM21_DATA20_SIG,
    DATA21 => ROM21_DATA21_SIG,
    DATA22 => ROM21_DATA22_SIG,
    DATA23 => ROM21_DATA23_SIG,
    DATA24 => ROM21_DATA24_SIG,
    DATA25 => ROM21_DATA25_SIG,
    DATA26 => ROM21_DATA26_SIG,
    DATA27 => ROM21_DATA27_SIG,
    DATA28 => ROM21_DATA28_SIG,
    DATA29 => ROM21_DATA29_SIG,
    DATA30 => ROM21_DATA30_SIG,
    DATA31 => ROM21_DATA31_SIG
);

WEIGHT_ROM22_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR22_0_SIG, 
    ADDR1  => ADDR22_1_SIG,
    ADDR2  => ADDR22_2_SIG,
    ADDR3  => ADDR22_3_SIG,
    ADDR4  => ADDR22_4_SIG,
    ADDR5  => ADDR22_5_SIG,
    ADDR6  => ADDR22_6_SIG,
    ADDR7  => ADDR22_7_SIG,
    ADDR8  => ADDR22_8_SIG,
    ADDR9  => ADDR22_9_SIG,
    ADDR10 => ADDR22_10_SIG,
    ADDR11 => ADDR22_11_SIG,
    ADDR12 => ADDR22_12_SIG,
    ADDR13 => ADDR22_13_SIG,
    ADDR14 => ADDR22_14_SIG,
    ADDR15 => ADDR22_15_SIG,
    ADDR16 => ADDR22_16_SIG,
    ADDR17 => ADDR22_17_SIG,
    ADDR18 => ADDR22_18_SIG,
    ADDR19 => ADDR22_19_SIG,
    ADDR20 => ADDR22_20_SIG,
    ADDR21 => ADDR22_21_SIG,
    ADDR22 => ADDR22_22_SIG,
    ADDR23 => ADDR22_23_SIG,
    ADDR24 => ADDR22_24_SIG,
    ADDR25 => ADDR22_25_SIG,
    ADDR26 => ADDR22_26_SIG,
    ADDR27 => ADDR22_27_SIG,
    ADDR28 => ADDR22_28_SIG,
    ADDR29 => ADDR22_29_SIG,
    ADDR30 => ADDR22_30_SIG,
    ADDR31 => ADDR22_31_SIG,
    DATA0  => ROM22_DATA0_SIG,
    DATA1  => ROM22_DATA1_SIG,
    DATA2  => ROM22_DATA2_SIG,
    DATA3  => ROM22_DATA3_SIG,
    DATA4  => ROM22_DATA4_SIG,
    DATA5  => ROM22_DATA5_SIG,
    DATA6  => ROM22_DATA6_SIG,
    DATA7  => ROM22_DATA7_SIG,
    DATA8  => ROM22_DATA8_SIG,
    DATA9  => ROM22_DATA9_SIG,
    DATA10 => ROM22_DATA10_SIG,
    DATA11 => ROM22_DATA11_SIG,
    DATA12 => ROM22_DATA12_SIG,
    DATA13 => ROM22_DATA13_SIG,
    DATA14 => ROM22_DATA14_SIG,
    DATA15 => ROM22_DATA15_SIG,
    DATA16 => ROM22_DATA16_SIG,
    DATA17 => ROM22_DATA17_SIG,
    DATA18 => ROM22_DATA18_SIG,
    DATA19 => ROM22_DATA19_SIG,
    DATA20 => ROM22_DATA20_SIG,
    DATA21 => ROM22_DATA21_SIG,
    DATA22 => ROM22_DATA22_SIG,
    DATA23 => ROM22_DATA23_SIG,
    DATA24 => ROM22_DATA24_SIG,
    DATA25 => ROM22_DATA25_SIG,
    DATA26 => ROM22_DATA26_SIG,
    DATA27 => ROM22_DATA27_SIG,
    DATA28 => ROM22_DATA28_SIG,
    DATA29 => ROM22_DATA29_SIG,
    DATA30 => ROM22_DATA30_SIG,
    DATA31 => ROM22_DATA31_SIG
);

WEIGHT_ROM23_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR23_0_SIG, 
    ADDR1  => ADDR23_1_SIG,
    ADDR2  => ADDR23_2_SIG,
    ADDR3  => ADDR23_3_SIG,
    ADDR4  => ADDR23_4_SIG,
    ADDR5  => ADDR23_5_SIG,
    ADDR6  => ADDR23_6_SIG,
    ADDR7  => ADDR23_7_SIG,
    ADDR8  => ADDR23_8_SIG,
    ADDR9  => ADDR23_9_SIG,
    ADDR10 => ADDR23_10_SIG,
    ADDR11 => ADDR23_11_SIG,
    ADDR12 => ADDR23_12_SIG,
    ADDR13 => ADDR23_13_SIG,
    ADDR14 => ADDR23_14_SIG,
    ADDR15 => ADDR23_15_SIG,
    ADDR16 => ADDR23_16_SIG,
    ADDR17 => ADDR23_17_SIG,
    ADDR18 => ADDR23_18_SIG,
    ADDR19 => ADDR23_19_SIG,
    ADDR20 => ADDR23_20_SIG,
    ADDR21 => ADDR23_21_SIG,
    ADDR22 => ADDR23_22_SIG,
    ADDR23 => ADDR23_23_SIG,
    ADDR24 => ADDR23_24_SIG,
    ADDR25 => ADDR23_25_SIG,
    ADDR26 => ADDR23_26_SIG,
    ADDR27 => ADDR23_27_SIG,
    ADDR28 => ADDR23_28_SIG,
    ADDR29 => ADDR23_29_SIG,
    ADDR30 => ADDR23_30_SIG,
    ADDR31 => ADDR23_31_SIG,
    DATA0  => ROM23_DATA0_SIG,
    DATA1  => ROM23_DATA1_SIG,
    DATA2  => ROM23_DATA2_SIG,
    DATA3  => ROM23_DATA3_SIG,
    DATA4  => ROM23_DATA4_SIG,
    DATA5  => ROM23_DATA5_SIG,
    DATA6  => ROM23_DATA6_SIG,
    DATA7  => ROM23_DATA7_SIG,
    DATA8  => ROM23_DATA8_SIG,
    DATA9  => ROM23_DATA9_SIG,
    DATA10 => ROM23_DATA10_SIG,
    DATA11 => ROM23_DATA11_SIG,
    DATA12 => ROM23_DATA12_SIG,
    DATA13 => ROM23_DATA13_SIG,
    DATA14 => ROM23_DATA14_SIG,
    DATA15 => ROM23_DATA15_SIG,
    DATA16 => ROM23_DATA16_SIG,
    DATA17 => ROM23_DATA17_SIG,
    DATA18 => ROM23_DATA18_SIG,
    DATA19 => ROM23_DATA19_SIG,
    DATA20 => ROM23_DATA20_SIG,
    DATA21 => ROM23_DATA21_SIG,
    DATA22 => ROM23_DATA22_SIG,
    DATA23 => ROM23_DATA23_SIG,
    DATA24 => ROM23_DATA24_SIG,
    DATA25 => ROM23_DATA25_SIG,
    DATA26 => ROM23_DATA26_SIG,
    DATA27 => ROM23_DATA27_SIG,
    DATA28 => ROM23_DATA28_SIG,
    DATA29 => ROM23_DATA29_SIG,
    DATA30 => ROM23_DATA30_SIG,
    DATA31 => ROM23_DATA31_SIG
);

WEIGHT_ROM24_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR24_0_SIG, 
    ADDR1  => ADDR24_1_SIG,
    ADDR2  => ADDR24_2_SIG,
    ADDR3  => ADDR24_3_SIG,
    ADDR4  => ADDR24_4_SIG,
    ADDR5  => ADDR24_5_SIG,
    ADDR6  => ADDR24_6_SIG,
    ADDR7  => ADDR24_7_SIG,
    ADDR8  => ADDR24_8_SIG,
    ADDR9  => ADDR24_9_SIG,
    ADDR10 => ADDR24_10_SIG,
    ADDR11 => ADDR24_11_SIG,
    ADDR12 => ADDR24_12_SIG,
    ADDR13 => ADDR24_13_SIG,
    ADDR14 => ADDR24_14_SIG,
    ADDR15 => ADDR24_15_SIG,
    ADDR16 => ADDR24_16_SIG,
    ADDR17 => ADDR24_17_SIG,
    ADDR18 => ADDR24_18_SIG,
    ADDR19 => ADDR24_19_SIG,
    ADDR20 => ADDR24_20_SIG,
    ADDR21 => ADDR24_21_SIG,
    ADDR22 => ADDR24_22_SIG,
    ADDR23 => ADDR24_23_SIG,
    ADDR24 => ADDR24_24_SIG,
    ADDR25 => ADDR24_25_SIG,
    ADDR26 => ADDR24_26_SIG,
    ADDR27 => ADDR24_27_SIG,
    ADDR28 => ADDR24_28_SIG,
    ADDR29 => ADDR24_29_SIG,
    ADDR30 => ADDR24_30_SIG,
    ADDR31 => ADDR24_31_SIG,
    DATA0  => ROM24_DATA0_SIG,
    DATA1  => ROM24_DATA1_SIG,
    DATA2  => ROM24_DATA2_SIG,
    DATA3  => ROM24_DATA3_SIG,
    DATA4  => ROM24_DATA4_SIG,
    DATA5  => ROM24_DATA5_SIG,
    DATA6  => ROM24_DATA6_SIG,
    DATA7  => ROM24_DATA7_SIG,
    DATA8  => ROM24_DATA8_SIG,
    DATA9  => ROM24_DATA9_SIG,
    DATA10 => ROM24_DATA10_SIG,
    DATA11 => ROM24_DATA11_SIG,
    DATA12 => ROM24_DATA12_SIG,
    DATA13 => ROM24_DATA13_SIG,
    DATA14 => ROM24_DATA14_SIG,
    DATA15 => ROM24_DATA15_SIG,
    DATA16 => ROM24_DATA16_SIG,
    DATA17 => ROM24_DATA17_SIG,
    DATA18 => ROM24_DATA18_SIG,
    DATA19 => ROM24_DATA19_SIG,
    DATA20 => ROM24_DATA20_SIG,
    DATA21 => ROM24_DATA21_SIG,
    DATA22 => ROM24_DATA22_SIG,
    DATA23 => ROM24_DATA23_SIG,
    DATA24 => ROM24_DATA24_SIG,
    DATA25 => ROM24_DATA25_SIG,
    DATA26 => ROM24_DATA26_SIG,
    DATA27 => ROM24_DATA27_SIG,
    DATA28 => ROM24_DATA28_SIG,
    DATA29 => ROM24_DATA29_SIG,
    DATA30 => ROM24_DATA30_SIG,
    DATA31 => ROM24_DATA31_SIG
);

WEIGHT_ROM25_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR25_0_SIG, 
    ADDR1  => ADDR25_1_SIG,
    ADDR2  => ADDR25_2_SIG,
    ADDR3  => ADDR25_3_SIG,
    ADDR4  => ADDR25_4_SIG,
    ADDR5  => ADDR25_5_SIG,
    ADDR6  => ADDR25_6_SIG,
    ADDR7  => ADDR25_7_SIG,
    ADDR8  => ADDR25_8_SIG,
    ADDR9  => ADDR25_9_SIG,
    ADDR10 => ADDR25_10_SIG,
    ADDR11 => ADDR25_11_SIG,
    ADDR12 => ADDR25_12_SIG,
    ADDR13 => ADDR25_13_SIG,
    ADDR14 => ADDR25_14_SIG,
    ADDR15 => ADDR25_15_SIG,
    ADDR16 => ADDR25_16_SIG,
    ADDR17 => ADDR25_17_SIG,
    ADDR18 => ADDR25_18_SIG,
    ADDR19 => ADDR25_19_SIG,
    ADDR20 => ADDR25_20_SIG,
    ADDR21 => ADDR25_21_SIG,
    ADDR22 => ADDR25_22_SIG,
    ADDR23 => ADDR25_23_SIG,
    ADDR24 => ADDR25_24_SIG,
    ADDR25 => ADDR25_25_SIG,
    ADDR26 => ADDR25_26_SIG,
    ADDR27 => ADDR25_27_SIG,
    ADDR28 => ADDR25_28_SIG,
    ADDR29 => ADDR25_29_SIG,
    ADDR30 => ADDR25_30_SIG,
    ADDR31 => ADDR25_31_SIG,
    DATA0  => ROM25_DATA0_SIG,
    DATA1  => ROM25_DATA1_SIG,
    DATA2  => ROM25_DATA2_SIG,
    DATA3  => ROM25_DATA3_SIG,
    DATA4  => ROM25_DATA4_SIG,
    DATA5  => ROM25_DATA5_SIG,
    DATA6  => ROM25_DATA6_SIG,
    DATA7  => ROM25_DATA7_SIG,
    DATA8  => ROM25_DATA8_SIG,
    DATA9  => ROM25_DATA9_SIG,
    DATA10 => ROM25_DATA10_SIG,
    DATA11 => ROM25_DATA11_SIG,
    DATA12 => ROM25_DATA12_SIG,
    DATA13 => ROM25_DATA13_SIG,
    DATA14 => ROM25_DATA14_SIG,
    DATA15 => ROM25_DATA15_SIG,
    DATA16 => ROM25_DATA16_SIG,
    DATA17 => ROM25_DATA17_SIG,
    DATA18 => ROM25_DATA18_SIG,
    DATA19 => ROM25_DATA19_SIG,
    DATA20 => ROM25_DATA20_SIG,
    DATA21 => ROM25_DATA21_SIG,
    DATA22 => ROM25_DATA22_SIG,
    DATA23 => ROM25_DATA23_SIG,
    DATA24 => ROM25_DATA24_SIG,
    DATA25 => ROM25_DATA25_SIG,
    DATA26 => ROM25_DATA26_SIG,
    DATA27 => ROM25_DATA27_SIG,
    DATA28 => ROM25_DATA28_SIG,
    DATA29 => ROM25_DATA29_SIG,
    DATA30 => ROM25_DATA30_SIG,
    DATA31 => ROM25_DATA31_SIG
);

WEIGHT_ROM26_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR26_0_SIG, 
    ADDR1  => ADDR26_1_SIG,
    ADDR2  => ADDR26_2_SIG,
    ADDR3  => ADDR26_3_SIG,
    ADDR4  => ADDR26_4_SIG,
    ADDR5  => ADDR26_5_SIG,
    ADDR6  => ADDR26_6_SIG,
    ADDR7  => ADDR26_7_SIG,
    ADDR8  => ADDR26_8_SIG,
    ADDR9  => ADDR26_9_SIG,
    ADDR10 => ADDR26_10_SIG,
    ADDR11 => ADDR26_11_SIG,
    ADDR12 => ADDR26_12_SIG,
    ADDR13 => ADDR26_13_SIG,
    ADDR14 => ADDR26_14_SIG,
    ADDR15 => ADDR26_15_SIG,
    ADDR16 => ADDR26_16_SIG,
    ADDR17 => ADDR26_17_SIG,
    ADDR18 => ADDR26_18_SIG,
    ADDR19 => ADDR26_19_SIG,
    ADDR20 => ADDR26_20_SIG,
    ADDR21 => ADDR26_21_SIG,
    ADDR22 => ADDR26_22_SIG,
    ADDR23 => ADDR26_23_SIG,
    ADDR24 => ADDR26_24_SIG,
    ADDR25 => ADDR26_25_SIG,
    ADDR26 => ADDR26_26_SIG,
    ADDR27 => ADDR26_27_SIG,
    ADDR28 => ADDR26_28_SIG,
    ADDR29 => ADDR26_29_SIG,
    ADDR30 => ADDR26_30_SIG,
    ADDR31 => ADDR26_31_SIG,
    DATA0  => ROM26_DATA0_SIG,
    DATA1  => ROM26_DATA1_SIG,
    DATA2  => ROM26_DATA2_SIG,
    DATA3  => ROM26_DATA3_SIG,
    DATA4  => ROM26_DATA4_SIG,
    DATA5  => ROM26_DATA5_SIG,
    DATA6  => ROM26_DATA6_SIG,
    DATA7  => ROM26_DATA7_SIG,
    DATA8  => ROM26_DATA8_SIG,
    DATA9  => ROM26_DATA9_SIG,
    DATA10 => ROM26_DATA10_SIG,
    DATA11 => ROM26_DATA11_SIG,
    DATA12 => ROM26_DATA12_SIG,
    DATA13 => ROM26_DATA13_SIG,
    DATA14 => ROM26_DATA14_SIG,
    DATA15 => ROM26_DATA15_SIG,
    DATA16 => ROM26_DATA16_SIG,
    DATA17 => ROM26_DATA17_SIG,
    DATA18 => ROM26_DATA18_SIG,
    DATA19 => ROM26_DATA19_SIG,
    DATA20 => ROM26_DATA20_SIG,
    DATA21 => ROM26_DATA21_SIG,
    DATA22 => ROM26_DATA22_SIG,
    DATA23 => ROM26_DATA23_SIG,
    DATA24 => ROM26_DATA24_SIG,
    DATA25 => ROM26_DATA25_SIG,
    DATA26 => ROM26_DATA26_SIG,
    DATA27 => ROM26_DATA27_SIG,
    DATA28 => ROM26_DATA28_SIG,
    DATA29 => ROM26_DATA29_SIG,
    DATA30 => ROM26_DATA30_SIG,
    DATA31 => ROM26_DATA31_SIG
);

WEIGHT_ROM27_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR27_0_SIG, 
    ADDR1  => ADDR27_1_SIG,
    ADDR2  => ADDR27_2_SIG,
    ADDR3  => ADDR27_3_SIG,
    ADDR4  => ADDR27_4_SIG,
    ADDR5  => ADDR27_5_SIG,
    ADDR6  => ADDR27_6_SIG,
    ADDR7  => ADDR27_7_SIG,
    ADDR8  => ADDR27_8_SIG,
    ADDR9  => ADDR27_9_SIG,
    ADDR10 => ADDR27_10_SIG,
    ADDR11 => ADDR27_11_SIG,
    ADDR12 => ADDR27_12_SIG,
    ADDR13 => ADDR27_13_SIG,
    ADDR14 => ADDR27_14_SIG,
    ADDR15 => ADDR27_15_SIG,
    ADDR16 => ADDR27_16_SIG,
    ADDR17 => ADDR27_17_SIG,
    ADDR18 => ADDR27_18_SIG,
    ADDR19 => ADDR27_19_SIG,
    ADDR20 => ADDR27_20_SIG,
    ADDR21 => ADDR27_21_SIG,
    ADDR22 => ADDR27_22_SIG,
    ADDR23 => ADDR27_23_SIG,
    ADDR24 => ADDR27_24_SIG,
    ADDR25 => ADDR27_25_SIG,
    ADDR26 => ADDR27_26_SIG,
    ADDR27 => ADDR27_27_SIG,
    ADDR28 => ADDR27_28_SIG,
    ADDR29 => ADDR27_29_SIG,
    ADDR30 => ADDR27_30_SIG,
    ADDR31 => ADDR27_31_SIG,
    DATA0  => ROM27_DATA0_SIG,
    DATA1  => ROM27_DATA1_SIG,
    DATA2  => ROM27_DATA2_SIG,
    DATA3  => ROM27_DATA3_SIG,
    DATA4  => ROM27_DATA4_SIG,
    DATA5  => ROM27_DATA5_SIG,
    DATA6  => ROM27_DATA6_SIG,
    DATA7  => ROM27_DATA7_SIG,
    DATA8  => ROM27_DATA8_SIG,
    DATA9  => ROM27_DATA9_SIG,
    DATA10 => ROM27_DATA10_SIG,
    DATA11 => ROM27_DATA11_SIG,
    DATA12 => ROM27_DATA12_SIG,
    DATA13 => ROM27_DATA13_SIG,
    DATA14 => ROM27_DATA14_SIG,
    DATA15 => ROM27_DATA15_SIG,
    DATA16 => ROM27_DATA16_SIG,
    DATA17 => ROM27_DATA17_SIG,
    DATA18 => ROM27_DATA18_SIG,
    DATA19 => ROM27_DATA19_SIG,
    DATA20 => ROM27_DATA20_SIG,
    DATA21 => ROM27_DATA21_SIG,
    DATA22 => ROM27_DATA22_SIG,
    DATA23 => ROM27_DATA23_SIG,
    DATA24 => ROM27_DATA24_SIG,
    DATA25 => ROM27_DATA25_SIG,
    DATA26 => ROM27_DATA26_SIG,
    DATA27 => ROM27_DATA27_SIG,
    DATA28 => ROM27_DATA28_SIG,
    DATA29 => ROM27_DATA29_SIG,
    DATA30 => ROM27_DATA30_SIG,
    DATA31 => ROM27_DATA31_SIG
);

WEIGHT_ROM28_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR28_0_SIG, 
    ADDR1  => ADDR28_1_SIG,
    ADDR2  => ADDR28_2_SIG,
    ADDR3  => ADDR28_3_SIG,
    ADDR4  => ADDR28_4_SIG,
    ADDR5  => ADDR28_5_SIG,
    ADDR6  => ADDR28_6_SIG,
    ADDR7  => ADDR28_7_SIG,
    ADDR8  => ADDR28_8_SIG,
    ADDR9  => ADDR28_9_SIG,
    ADDR10 => ADDR28_10_SIG,
    ADDR11 => ADDR28_11_SIG,
    ADDR12 => ADDR28_12_SIG,
    ADDR13 => ADDR28_13_SIG,
    ADDR14 => ADDR28_14_SIG,
    ADDR15 => ADDR28_15_SIG,
    ADDR16 => ADDR28_16_SIG,
    ADDR17 => ADDR28_17_SIG,
    ADDR18 => ADDR28_18_SIG,
    ADDR19 => ADDR28_19_SIG,
    ADDR20 => ADDR28_20_SIG,
    ADDR21 => ADDR28_21_SIG,
    ADDR22 => ADDR28_22_SIG,
    ADDR23 => ADDR28_23_SIG,
    ADDR24 => ADDR28_24_SIG,
    ADDR25 => ADDR28_25_SIG,
    ADDR26 => ADDR28_26_SIG,
    ADDR27 => ADDR28_27_SIG,
    ADDR28 => ADDR28_28_SIG,
    ADDR29 => ADDR28_29_SIG,
    ADDR30 => ADDR28_30_SIG,
    ADDR31 => ADDR28_31_SIG,
    DATA0  => ROM28_DATA0_SIG,
    DATA1  => ROM28_DATA1_SIG,
    DATA2  => ROM28_DATA2_SIG,
    DATA3  => ROM28_DATA3_SIG,
    DATA4  => ROM28_DATA4_SIG,
    DATA5  => ROM28_DATA5_SIG,
    DATA6  => ROM28_DATA6_SIG,
    DATA7  => ROM28_DATA7_SIG,
    DATA8  => ROM28_DATA8_SIG,
    DATA9  => ROM28_DATA9_SIG,
    DATA10 => ROM28_DATA10_SIG,
    DATA11 => ROM28_DATA11_SIG,
    DATA12 => ROM28_DATA12_SIG,
    DATA13 => ROM28_DATA13_SIG,
    DATA14 => ROM28_DATA14_SIG,
    DATA15 => ROM28_DATA15_SIG,
    DATA16 => ROM28_DATA16_SIG,
    DATA17 => ROM28_DATA17_SIG,
    DATA18 => ROM28_DATA18_SIG,
    DATA19 => ROM28_DATA19_SIG,
    DATA20 => ROM28_DATA20_SIG,
    DATA21 => ROM28_DATA21_SIG,
    DATA22 => ROM28_DATA22_SIG,
    DATA23 => ROM28_DATA23_SIG,
    DATA24 => ROM28_DATA24_SIG,
    DATA25 => ROM28_DATA25_SIG,
    DATA26 => ROM28_DATA26_SIG,
    DATA27 => ROM28_DATA27_SIG,
    DATA28 => ROM28_DATA28_SIG,
    DATA29 => ROM28_DATA29_SIG,
    DATA30 => ROM28_DATA30_SIG,
    DATA31 => ROM28_DATA31_SIG
);

WEIGHT_ROM29_INST: WEIGHT_ROM
Generic map ( WIDTH => 32, POWER => 13)
Port map(
    ADDR0  => ADDR29_0_SIG, 
    ADDR1  => ADDR29_1_SIG,
    ADDR2  => ADDR29_2_SIG,
    ADDR3  => ADDR29_3_SIG,
    ADDR4  => ADDR29_4_SIG,
    ADDR5  => ADDR29_5_SIG,
    ADDR6  => ADDR29_6_SIG,
    ADDR7  => ADDR29_7_SIG,
    ADDR8  => ADDR29_8_SIG,
    ADDR9  => ADDR29_9_SIG,
    ADDR10 => ADDR29_10_SIG,
    ADDR11 => ADDR29_11_SIG,
    ADDR12 => ADDR29_12_SIG,
    ADDR13 => ADDR29_13_SIG,
    ADDR14 => ADDR29_14_SIG,
    ADDR15 => ADDR29_15_SIG,
    ADDR16 => ADDR29_16_SIG,
    ADDR17 => ADDR29_17_SIG,
    ADDR18 => ADDR29_18_SIG,
    ADDR19 => ADDR29_19_SIG,
    ADDR20 => ADDR29_20_SIG,
    ADDR21 => ADDR29_21_SIG,
    ADDR22 => ADDR29_22_SIG,
    ADDR23 => ADDR29_23_SIG,
    ADDR24 => ADDR29_24_SIG,
    ADDR25 => ADDR29_25_SIG,
    ADDR26 => ADDR29_26_SIG,
    ADDR27 => ADDR29_27_SIG,
    ADDR28 => ADDR29_28_SIG,
    ADDR29 => ADDR29_29_SIG,
    ADDR30 => ADDR29_30_SIG,
    ADDR31 => ADDR29_31_SIG,
    DATA0  => ROM29_DATA0_SIG,
    DATA1  => ROM29_DATA1_SIG,
    DATA2  => ROM29_DATA2_SIG,
    DATA3  => ROM29_DATA3_SIG,
    DATA4  => ROM29_DATA4_SIG,
    DATA5  => ROM29_DATA5_SIG,
    DATA6  => ROM29_DATA6_SIG,
    DATA7  => ROM29_DATA7_SIG,
    DATA8  => ROM29_DATA8_SIG,
    DATA9  => ROM29_DATA9_SIG,
    DATA10 => ROM29_DATA10_SIG,
    DATA11 => ROM29_DATA11_SIG,
    DATA12 => ROM29_DATA12_SIG,
    DATA13 => ROM29_DATA13_SIG,
    DATA14 => ROM29_DATA14_SIG,
    DATA15 => ROM29_DATA15_SIG,
    DATA16 => ROM29_DATA16_SIG,
    DATA17 => ROM29_DATA17_SIG,
    DATA18 => ROM29_DATA18_SIG,
    DATA19 => ROM29_DATA19_SIG,
    DATA20 => ROM29_DATA20_SIG,
    DATA21 => ROM29_DATA21_SIG,
    DATA22 => ROM29_DATA22_SIG,
    DATA23 => ROM29_DATA23_SIG,
    DATA24 => ROM29_DATA24_SIG,
    DATA25 => ROM29_DATA25_SIG,
    DATA26 => ROM29_DATA26_SIG,
    DATA27 => ROM29_DATA27_SIG,
    DATA28 => ROM29_DATA28_SIG,
    DATA29 => ROM29_DATA29_SIG,
    DATA30 => ROM29_DATA30_SIG,
    DATA31 => ROM29_DATA31_SIG
);

BIAS_ROM_INST: BIAS_ROM_FC
Generic map ( WIDTH => 64, POWER => 5 )
Port map (
    ADDR0  => BIAS0_ROM_ADDR,
    ADDR1  => BIAS1_ROM_ADDR, 
    ADDR2  => BIAS2_ROM_ADDR,
    ADDR3  => BIAS3_ROM_ADDR,
    ADDR4  => BIAS4_ROM_ADDR,
    ADDR5  => BIAS5_ROM_ADDR,
    ADDR6  => BIAS6_ROM_ADDR,
    ADDR7  => BIAS7_ROM_ADDR,
    ADDR8  => BIAS8_ROM_ADDR,
    ADDR9  => BIAS9_ROM_ADDR,
    ADDR10 => BIAS10_ROM_ADDR,
    ADDR11 => BIAS11_ROM_ADDR,
    ADDR12 => BIAS12_ROM_ADDR,
    ADDR13 => BIAS13_ROM_ADDR,
    ADDR14 => BIAS14_ROM_ADDR,
    ADDR15 => BIAS15_ROM_ADDR,
    ADDR16 => BIAS16_ROM_ADDR,
    ADDR17 => BIAS17_ROM_ADDR,
    ADDR18 => BIAS18_ROM_ADDR,
    ADDR19 => BIAS19_ROM_ADDR,
    ADDR20 => BIAS20_ROM_ADDR,
    ADDR21 => BIAS21_ROM_ADDR,
    ADDR22 => BIAS22_ROM_ADDR,
    ADDR23 => BIAS23_ROM_ADDR,
    ADDR24 => BIAS24_ROM_ADDR,
    ADDR25 => BIAS25_ROM_ADDR,
    ADDR26 => BIAS26_ROM_ADDR,
    ADDR27 => BIAS27_ROM_ADDR,
    ADDR28 => BIAS28_ROM_ADDR,
    ADDR29 => BIAS29_ROM_ADDR,
    DATA0  => BIAS0_SIG,
    DATA1  => BIAS1_SIG,
    DATA2  => BIAS2_SIG,
    DATA3  => BIAS3_SIG,
    DATA4  => BIAS4_SIG,
    DATA5  => BIAS5_SIG,
    DATA6  => BIAS6_SIG,
    DATA7  => BIAS7_SIG,
    DATA8  => BIAS8_SIG,
    DATA9  => BIAS9_SIG,
    DATA10 => BIAS10_SIG,
    DATA11 => BIAS11_SIG,
    DATA12 => BIAS12_SIG,
    DATA13 => BIAS13_SIG,
    DATA14 => BIAS14_SIG,
    DATA15 => BIAS15_SIG,
    DATA16 => BIAS16_SIG,
    DATA17 => BIAS17_SIG,
    DATA18 => BIAS18_SIG,
    DATA19 => BIAS19_SIG,
    DATA20 => BIAS20_SIG,
    DATA21 => BIAS21_SIG,
    DATA22 => BIAS22_SIG,
    DATA23 => BIAS23_SIG,
    DATA24 => BIAS24_SIG,
    DATA25 => BIAS25_SIG,
    DATA26 => BIAS26_SIG,
    DATA27 => BIAS27_SIG,
    DATA28 => BIAS28_SIG,
    DATA29 => BIAS29_SIG
);

ADDER0_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS0_SIG,
    B    => VM0_OUT_SIG,
    S    => ADDER0_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER1_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS1_SIG,
    B    => VM1_OUT_SIG,
    S    => ADDER1_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER2_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS2_SIG,
    B    => VM2_OUT_SIG,
    S    => ADDER2_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER3_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS3_SIG,
    B    => VM3_OUT_SIG,
    S    => ADDER3_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER4_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS4_SIG,
    B    => VM4_OUT_SIG,
    S    => ADDER4_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER5_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS5_SIG,
    B    => VM5_OUT_SIG,
    S    => ADDER5_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER6_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS6_SIG,
    B    => VM6_OUT_SIG,
    S    => ADDER6_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER7_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS7_SIG,
    B    => VM7_OUT_SIG,
    S    => ADDER7_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER8_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS8_SIG,
    B    => VM8_OUT_SIG,
    S    => ADDER8_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER9_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS9_SIG,
    B    => VM9_OUT_SIG,
    S    => ADDER9_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER10_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS10_SIG,
    B    => VM10_OUT_SIG,
    S    => ADDER10_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER11_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS11_SIG,
    B    => VM11_OUT_SIG,
    S    => ADDER11_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER12_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS12_SIG,
    B    => VM12_OUT_SIG,
    S    => ADDER12_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER13_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS13_SIG,
    B    => VM13_OUT_SIG,
    S    => ADDER13_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER14_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS14_SIG,
    B    => VM14_OUT_SIG,
    S    => ADDER14_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER15_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS15_SIG,
    B    => VM15_OUT_SIG,
    S    => ADDER15_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER16_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS16_SIG,
    B    => VM16_OUT_SIG,
    S    => ADDER16_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER17_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS17_SIG,
    B    => VM17_OUT_SIG,
    S    => ADDER17_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER18_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS18_SIG,
    B    => VM18_OUT_SIG,
    S    => ADDER18_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER19_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS19_SIG,
    B    => VM19_OUT_SIG,
    S    => ADDER19_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER20_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS20_SIG,
    B    => VM20_OUT_SIG,
    S    => ADDER20_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER21_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS21_SIG,
    B    => VM21_OUT_SIG,
    S    => ADDER21_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER22_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS22_SIG,
    B    => VM22_OUT_SIG,
    S    => ADDER22_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER23_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS23_SIG,
    B    => VM23_OUT_SIG,
    S    => ADDER23_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER24_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS24_SIG,
    B    => VM24_OUT_SIG,
    S    => ADDER24_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER25_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS25_SIG,
    B    => VM25_OUT_SIG,
    S    => ADDER25_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER26_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS26_SIG,
    B    => VM26_OUT_SIG,
    S    => ADDER26_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER27_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS27_SIG,
    B    => VM27_OUT_SIG,
    S    => ADDER27_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER28_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS28_SIG,
    B    => VM28_OUT_SIG,
    S    => ADDER28_OUT_SIG,
    COUT => open,
    OV   => open
);

ADDER29_INST: ADDER
Generic map ( WIDTH => 64)
Port map (
    A    => BIAS29_SIG,
    B    => VM29_OUT_SIG,
    S    => ADDER29_OUT_SIG,
    COUT => open,
    OV   => open
);

RELU_MUX0_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER0_OUT_SIG,
    DOUT  => DOUT0
);

RELU_MUX1_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER1_OUT_SIG,
    DOUT  => DOUT1
);

RELU_MUX2_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER2_OUT_SIG,
    DOUT  => DOUT2
);

RELU_MUX3_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER3_OUT_SIG,
    DOUT  => DOUT3
);

RELU_MUX4_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER4_OUT_SIG,
    DOUT  => DOUT4
);

RELU_MUX5_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER5_OUT_SIG,
    DOUT  => DOUT5
);

RELU_MUX6_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER6_OUT_SIG,
    DOUT  => DOUT6
);

RELU_MUX7_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER7_OUT_SIG,
    DOUT  => DOUT7
);

RELU_MUX8_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER8_OUT_SIG,
    DOUT  => DOUT8
);

RELU_MUX9_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER9_OUT_SIG,
    DOUT  => DOUT9
);

RELU_MUX10_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER10_OUT_SIG,
    DOUT  => DOUT10
);

RELU_MUX11_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER11_OUT_SIG,
    DOUT  => DOUT11
);

RELU_MUX12_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER12_OUT_SIG,
    DOUT  => DOUT12
);

RELU_MUX13_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER13_OUT_SIG,
    DOUT  => DOUT13
);

RELU_MUX14_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER14_OUT_SIG,
    DOUT  => DOUT14
);

RELU_MUX15_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER15_OUT_SIG,
    DOUT  => DOUT15
);

RELU_MUX16_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER16_OUT_SIG,
    DOUT  => DOUT16
);

RELU_MUX17_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER17_OUT_SIG,
    DOUT  => DOUT17
);

RELU_MUX18_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER18_OUT_SIG,
    DOUT  => DOUT18
);

RELU_MUX19_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER19_OUT_SIG,
    DOUT  => DOUT19
);

RELU_MUX20_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER20_OUT_SIG,
    DOUT  => DOUT20
);

RELU_MUX21_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER21_OUT_SIG,
    DOUT  => DOUT21
);

RELU_MUX22_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER22_OUT_SIG,
    DOUT  => DOUT22
);

RELU_MUX23_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER23_OUT_SIG,
    DOUT  => DOUT23
);

RELU_MUX24_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER24_OUT_SIG,
    DOUT  => DOUT24
);

RELU_MUX25_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER25_OUT_SIG,
    DOUT  => DOUT25
);

RELU_MUX26_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER26_OUT_SIG,
    DOUT  => DOUT26
);

RELU_MUX27_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER27_OUT_SIG,
    DOUT  => DOUT27
);

RELU_MUX28_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER28_OUT_SIG,
    DOUT  => DOUT28
);

RELU_MUX29_INST: RELU_MUX
Generic map ( WIDTH => 64 )
Port map (
    DIN   => ADDER29_OUT_SIG,
    DOUT  => DOUT29
);

end Structural;
