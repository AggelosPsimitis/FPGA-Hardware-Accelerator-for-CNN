library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity CONVOLUTION_LAYER is
Generic ( WIDTH : positive := 16);
Port (
    CLK    :  in   std_logic;
    RESET  :  in   std_logic;
    DIN0   :  in   std_logic_vector(WIDTH-1 downto 0);
    DIN1   :  in   std_logic_vector(WIDTH-1 downto 0);
    DIN2   :  in   std_logic_vector(WIDTH-1 downto 0);
    DIN3   :  in   std_logic_vector(WIDTH-1 downto 0);
    DIN4   :  in   std_logic_vector(WIDTH-1 downto 0);
    DOUT0  :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT1  :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT2  :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT3  :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT4  :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT5  :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT6  :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT7  :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT8  :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT9  :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT10 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT11 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT12 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT13 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT14 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT15 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT16 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT17 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT18 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT19 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT20 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT21 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT22 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT23 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT24 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT25 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT26 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT27 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT28 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT29 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT30 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0);
    DOUT31 :  out  std_logic_vector(WIDTH+WIDTH-1 downto 0)
);
end CONVOLUTION_LAYER;

architecture Structural of CONVOLUTION_LAYER is

component DSP_BLOCK
Generic ( PIXEL_SIZE : positive := 16;
          POWER : positive := 5);
Port (
    CLK       :  in  std_logic;
    RESET     :  in  std_logic;
    DIN0      :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    DIN1      :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    DIN2      :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    DIN3      :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    DIN4      :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE00_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE01_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE02_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE03_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE04_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE10_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE11_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE12_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE13_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE14_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE20_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE21_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE22_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE23_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE24_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE30_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE31_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE32_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE33_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE34_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE40_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE41_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE42_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE43_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    PE44_COEF :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    BIAS      :  in  std_logic_vector(PIXEL_SIZE-1 downto 0);
    DOUT      :  out std_logic_vector(PIXEL_SIZE+PIXEL_SIZE-1 downto 0)
);
end component;

component ROM0 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM1 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM2 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM3 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM4 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM5 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM6 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM7 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM8 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM9 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM10 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM11 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM12 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM13 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM14 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM15 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM16 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM17 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM18 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM19 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM20 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM21 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM22 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM23 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM24 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM25 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM26 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM27
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM28 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM29 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM30 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

component ROM31 
Generic ( WIDTH : positive := 16;
          POWER : positive := 5); 
Port ( 
    ADDR0  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR1  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR2  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR3  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR4  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR5  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR6  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR7  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR8  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR9  :    in  std_logic_vector(POWER-1 downto 0);
    ADDR10 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR11 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR12 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR13 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR14 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR15 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR16 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR17 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR18 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR19 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR20 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR21 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR22 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR23 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR24 :    in  std_logic_vector(POWER-1 downto 0);
    ADDR25 :    in  std_logic_vector(POWER-1 downto 0);
    DATA0  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA1  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA2  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA3  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA4  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA5  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA6  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA7  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA8  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA9  :    out std_logic_vector(WIDTH-1 downto 0);
    DATA10 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA11 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA12 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA13 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA14 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA15 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA16 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA17 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA18 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA19 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA20 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA21 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA22 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA23 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA24 :    out std_logic_vector(WIDTH-1 downto 0);
    DATA25 :    out std_logic_vector(WIDTh-1 downto 0)
);
end component;

signal DIN0_SIG, DIN1_SIG, DIN2_SIG, DIN3_SIG, DIN4_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal DOUT0_SIG, DOUT1_SIG, DOUT2_SIG, DOUT3_SIG, DOUT4_SIG,
       DOUT5_SIG, DOUT6_SIG, DOUT7_SIG, DOUT8_SIG, DOUT9_SIG,
       DOUT10_SIG, DOUT11_SIG, DOUT12_SIG, DOUT13_SIG, DOUT14_SIG,
       DOUT15_SIG, DOUT16_SIG, DOUT17_SIG, DOUT18_SIG, DOUT19_SIG,
       DOUT20_SIG, DOUT21_SIG, DOUT22_SIG, DOUT23_SIG, DOUT24_SIG,
       DOUT25_SIG, DOUT26_SIG, DOUT27_SIG, DOUT28_SIG, DOUT29_SIG, DOUT30_SIG, DOUT31_SIG : std_logic_vector(WIDTH+WIDTH-1 downto 0) := (others => '0');
signal ADDR0_SIG  : std_logic_vector(4 downto 0) := "00000";
signal ADDR1_SIG  : std_logic_vector(4 downto 0) := "00001";
signal ADDR2_SIG  : std_logic_vector(4 downto 0) := "00010";
signal ADDR3_SIG  : std_logic_vector(4 downto 0) := "00011";
signal ADDR4_SIG  : std_logic_vector(4 downto 0) := "00100";
signal ADDR5_SIG  : std_logic_vector(4 downto 0) := "00101";
signal ADDR6_SIG  : std_logic_vector(4 downto 0) := "00110";
signal ADDR7_SIG  : std_logic_vector(4 downto 0) := "00111";
signal ADDR8_SIG  : std_logic_vector(4 downto 0) := "01000";
signal ADDR9_SIG  : std_logic_vector(4 downto 0) := "01001";
signal ADDR10_SIG : std_logic_vector(4 downto 0) := "01010";
signal ADDR11_SIG : std_logic_vector(4 downto 0) := "01011";
signal ADDR12_SIG : std_logic_vector(4 downto 0) := "01100";
signal ADDR13_SIG : std_logic_vector(4 downto 0) := "01101";
signal ADDR14_SIG : std_logic_vector(4 downto 0) := "01110";
signal ADDR15_SIG : std_logic_vector(4 downto 0) := "01111";
signal ADDR16_SIG : std_logic_vector(4 downto 0) := "10000";
signal ADDR17_SIG : std_logic_vector(4 downto 0) := "10001";
signal ADDR18_SIG : std_logic_vector(4 downto 0) := "10010";
signal ADDR19_SIG : std_logic_vector(4 downto 0) := "10011";
signal ADDR20_SIG : std_logic_vector(4 downto 0) := "10100";
signal ADDR21_SIG : std_logic_vector(4 downto 0) := "10101";
signal ADDR22_SIG : std_logic_vector(4 downto 0) := "10110";
signal ADDR23_SIG : std_logic_vector(4 downto 0) := "10111";
signal ADDR24_SIG : std_logic_vector(4 downto 0) := "11000";
signal ADDR25_SIG : std_logic_vector(4 downto 0) := "11001";
signal ROM0_DATA0_SIG, ROM0_DATA1_SIG, ROM0_DATA2_SIG, ROM0_DATA3_SIG, ROM0_DATA4_SIG,
       ROM0_DATA5_SIG, ROM0_DATA6_SIG, ROM0_DATA7_SIG, ROM0_DATA8_SIG, ROM0_DATA9_SIG,
       ROM0_DATA10_SIG, ROM0_DATA11_SIG, ROM0_DATA12_SIG, ROM0_DATA13_SIG, ROM0_DATA14_SIG,
       ROM0_DATA15_SIG, ROM0_DATA16_SIG, ROM0_DATA17_SIG, ROM0_DATA18_SIG, ROM0_DATA19_SIG,
       ROM0_DATA20_SIG, ROM0_DATA21_SIG, ROM0_DATA22_SIG, ROM0_DATA23_SIG, ROM0_DATA24_SIG, ROM0_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM1_DATA0_SIG, ROM1_DATA1_SIG, ROM1_DATA2_SIG, ROM1_DATA3_SIG, ROM1_DATA4_SIG,
       ROM1_DATA5_SIG, ROM1_DATA6_SIG, ROM1_DATA7_SIG, ROM1_DATA8_SIG, ROM1_DATA9_SIG,
       ROM1_DATA10_SIG, ROM1_DATA11_SIG, ROM1_DATA12_SIG, ROM1_DATA13_SIG, ROM1_DATA14_SIG,
       ROM1_DATA15_SIG, ROM1_DATA16_SIG, ROM1_DATA17_SIG, ROM1_DATA18_SIG, ROM1_DATA19_SIG,
       ROM1_DATA20_SIG, ROM1_DATA21_SIG, ROM1_DATA22_SIG, ROM1_DATA23_SIG, ROM1_DATA24_SIG, ROM1_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0'); 
signal ROM2_DATA0_SIG, ROM2_DATA1_SIG, ROM2_DATA2_SIG, ROM2_DATA3_SIG, ROM2_DATA4_SIG,
       ROM2_DATA5_SIG, ROM2_DATA6_SIG, ROM2_DATA7_SIG, ROM2_DATA8_SIG, ROM2_DATA9_SIG,
       ROM2_DATA10_SIG, ROM2_DATA11_SIG, ROM2_DATA12_SIG, ROM2_DATA13_SIG, ROM2_DATA14_SIG,
       ROM2_DATA15_SIG, ROM2_DATA16_SIG, ROM2_DATA17_SIG, ROM2_DATA18_SIG, ROM2_DATA19_SIG,
       ROM2_DATA20_SIG, ROM2_DATA21_SIG, ROM2_DATA22_SIG, ROM2_DATA23_SIG, ROM2_DATA24_SIG, ROM2_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM3_DATA0_SIG, ROM3_DATA1_SIG, ROM3_DATA2_SIG, ROM3_DATA3_SIG, ROM3_DATA4_SIG,
       ROM3_DATA5_SIG, ROM3_DATA6_SIG, ROM3_DATA7_SIG, ROM3_DATA8_SIG, ROM3_DATA9_SIG,
       ROM3_DATA10_SIG, ROM3_DATA11_SIG, ROM3_DATA12_SIG, ROM3_DATA13_SIG, ROM3_DATA14_SIG,
       ROM3_DATA15_SIG, ROM3_DATA16_SIG, ROM3_DATA17_SIG, ROM3_DATA18_SIG, ROM3_DATA19_SIG,
       ROM3_DATA20_SIG, ROM3_DATA21_SIG, ROM3_DATA22_SIG, ROM3_DATA23_SIG, ROM3_DATA24_SIG, ROM3_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM4_DATA0_SIG, ROM4_DATA1_SIG, ROM4_DATA2_SIG, ROM4_DATA3_SIG, ROM4_DATA4_SIG,
       ROM4_DATA5_SIG, ROM4_DATA6_SIG, ROM4_DATA7_SIG, ROM4_DATA8_SIG, ROM4_DATA9_SIG,
       ROM4_DATA10_SIG, ROM4_DATA11_SIG, ROM4_DATA12_SIG, ROM4_DATA13_SIG, ROM4_DATA14_SIG,
       ROM4_DATA15_SIG, ROM4_DATA16_SIG, ROM4_DATA17_SIG, ROM4_DATA18_SIG, ROM4_DATA19_SIG,
       ROM4_DATA20_SIG, ROM4_DATA21_SIG, ROM4_DATA22_SIG, ROM4_DATA23_SIG, ROM4_DATA24_SIG, ROM4_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0'); 
signal ROM5_DATA0_SIG, ROM5_DATA1_SIG, ROM5_DATA2_SIG, ROM5_DATA3_SIG, ROM5_DATA4_SIG,
       ROM5_DATA5_SIG, ROM5_DATA6_SIG, ROM5_DATA7_SIG, ROM5_DATA8_SIG, ROM5_DATA9_SIG,
       ROM5_DATA10_SIG, ROM5_DATA11_SIG, ROM5_DATA12_SIG, ROM5_DATA13_SIG, ROM5_DATA14_SIG,
       ROM5_DATA15_SIG, ROM5_DATA16_SIG, ROM5_DATA17_SIG, ROM5_DATA18_SIG, ROM5_DATA19_SIG,
       ROM5_DATA20_SIG, ROM5_DATA21_SIG, ROM5_DATA22_SIG, ROM5_DATA23_SIG, ROM5_DATA24_SIG, ROM5_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM6_DATA0_SIG, ROM6_DATA1_SIG, ROM6_DATA2_SIG, ROM6_DATA3_SIG, ROM6_DATA4_SIG,
       ROM6_DATA5_SIG, ROM6_DATA6_SIG, ROM6_DATA7_SIG, ROM6_DATA8_SIG, ROM6_DATA9_SIG,
       ROM6_DATA10_SIG, ROM6_DATA11_SIG, ROM6_DATA12_SIG, ROM6_DATA13_SIG, ROM6_DATA14_SIG,
       ROM6_DATA15_SIG, ROM6_DATA16_SIG, ROM6_DATA17_SIG, ROM6_DATA18_SIG, ROM6_DATA19_SIG,
       ROM6_DATA20_SIG, ROM6_DATA21_SIG, ROM6_DATA22_SIG, ROM6_DATA23_SIG, ROM6_DATA24_SIG, ROM6_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');   
signal ROM7_DATA0_SIG, ROM7_DATA1_SIG, ROM7_DATA2_SIG, ROM7_DATA3_SIG, ROM7_DATA4_SIG,
       ROM7_DATA5_SIG, ROM7_DATA6_SIG, ROM7_DATA7_SIG, ROM7_DATA8_SIG, ROM7_DATA9_SIG,
       ROM7_DATA10_SIG, ROM7_DATA11_SIG, ROM7_DATA12_SIG, ROM7_DATA13_SIG, ROM7_DATA14_SIG,
       ROM7_DATA15_SIG, ROM7_DATA16_SIG, ROM7_DATA17_SIG, ROM7_DATA18_SIG, ROM7_DATA19_SIG,
       ROM7_DATA20_SIG, ROM7_DATA21_SIG, ROM7_DATA22_SIG, ROM7_DATA23_SIG, ROM7_DATA24_SIG, ROM7_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0'); 
signal ROM8_DATA0_SIG, ROM8_DATA1_SIG, ROM8_DATA2_SIG, ROM8_DATA3_SIG, ROM8_DATA4_SIG,
       ROM8_DATA5_SIG, ROM8_DATA6_SIG, ROM8_DATA7_SIG, ROM8_DATA8_SIG, ROM8_DATA9_SIG,
       ROM8_DATA10_SIG, ROM8_DATA11_SIG, ROM8_DATA12_SIG, ROM8_DATA13_SIG, ROM8_DATA14_SIG,
       ROM8_DATA15_SIG, ROM8_DATA16_SIG, ROM8_DATA17_SIG, ROM8_DATA18_SIG, ROM8_DATA19_SIG,
       ROM8_DATA20_SIG, ROM8_DATA21_SIG, ROM8_DATA22_SIG, ROM8_DATA23_SIG, ROM8_DATA24_SIG, ROM8_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0'); 
signal ROM9_DATA0_SIG, ROM9_DATA1_SIG, ROM9_DATA2_SIG, ROM9_DATA3_SIG, ROM9_DATA4_SIG,
       ROM9_DATA5_SIG, ROM9_DATA6_SIG, ROM9_DATA7_SIG, ROM9_DATA8_SIG, ROM9_DATA9_SIG,
       ROM9_DATA10_SIG, ROM9_DATA11_SIG, ROM9_DATA12_SIG, ROM9_DATA13_SIG, ROM9_DATA14_SIG,
       ROM9_DATA15_SIG, ROM9_DATA16_SIG, ROM9_DATA17_SIG, ROM9_DATA18_SIG, ROM9_DATA19_SIG,
       ROM9_DATA20_SIG, ROM9_DATA21_SIG, ROM9_DATA22_SIG, ROM9_DATA23_SIG, ROM9_DATA24_SIG, ROM9_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0'); 
signal ROM10_DATA0_SIG, ROM10_DATA1_SIG, ROM10_DATA2_SIG, ROM10_DATA3_SIG, ROM10_DATA4_SIG,
       ROM10_DATA5_SIG, ROM10_DATA6_SIG, ROM10_DATA7_SIG, ROM10_DATA8_SIG, ROM10_DATA9_SIG,
       ROM10_DATA10_SIG, ROM10_DATA11_SIG, ROM10_DATA12_SIG, ROM10_DATA13_SIG, ROM10_DATA14_SIG,
       ROM10_DATA15_SIG, ROM10_DATA16_SIG, ROM10_DATA17_SIG, ROM10_DATA18_SIG, ROM10_DATA19_SIG,
       ROM10_DATA20_SIG, ROM10_DATA21_SIG, ROM10_DATA22_SIG, ROM10_DATA23_SIG, ROM10_DATA24_SIG, ROM10_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0'); 
signal ROM11_DATA0_SIG, ROM11_DATA1_SIG, ROM11_DATA2_SIG, ROM11_DATA3_SIG, ROM11_DATA4_SIG,
       ROM11_DATA5_SIG, ROM11_DATA6_SIG, ROM11_DATA7_SIG, ROM11_DATA8_SIG, ROM11_DATA9_SIG,
       ROM11_DATA10_SIG, ROM11_DATA11_SIG, ROM11_DATA12_SIG, ROM11_DATA13_SIG, ROM11_DATA14_SIG,
       ROM11_DATA15_SIG, ROM11_DATA16_SIG, ROM11_DATA17_SIG, ROM11_DATA18_SIG, ROM11_DATA19_SIG,
       ROM11_DATA20_SIG, ROM11_DATA21_SIG, ROM11_DATA22_SIG, ROM11_DATA23_SIG, ROM11_DATA24_SIG, ROM11_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0'); 
signal ROM12_DATA0_SIG, ROM12_DATA1_SIG, ROM12_DATA2_SIG, ROM12_DATA3_SIG, ROM12_DATA4_SIG,
       ROM12_DATA5_SIG, ROM12_DATA6_SIG, ROM12_DATA7_SIG, ROM12_DATA8_SIG, ROM12_DATA9_SIG,
       ROM12_DATA10_SIG, ROM12_DATA11_SIG, ROM12_DATA12_SIG, ROM12_DATA13_SIG, ROM12_DATA14_SIG,
       ROM12_DATA15_SIG, ROM12_DATA16_SIG, ROM12_DATA17_SIG, ROM12_DATA18_SIG, ROM12_DATA19_SIG,
       ROM12_DATA20_SIG, ROM12_DATA21_SIG, ROM12_DATA22_SIG, ROM12_DATA23_SIG, ROM12_DATA24_SIG, ROM12_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0'); 
signal ROM13_DATA0_SIG, ROM13_DATA1_SIG, ROM13_DATA2_SIG, ROM13_DATA3_SIG, ROM13_DATA4_SIG,
       ROM13_DATA5_SIG, ROM13_DATA6_SIG, ROM13_DATA7_SIG, ROM13_DATA8_SIG, ROM13_DATA9_SIG,
       ROM13_DATA10_SIG, ROM13_DATA11_SIG, ROM13_DATA12_SIG, ROM13_DATA13_SIG, ROM13_DATA14_SIG,
       ROM13_DATA15_SIG, ROM13_DATA16_SIG, ROM13_DATA17_SIG, ROM13_DATA18_SIG, ROM13_DATA19_SIG,
       ROM13_DATA20_SIG, ROM13_DATA21_SIG, ROM13_DATA22_SIG, ROM13_DATA23_SIG, ROM13_DATA24_SIG, ROM13_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0'); 
signal ROM14_DATA0_SIG, ROM14_DATA1_SIG, ROM14_DATA2_SIG, ROM14_DATA3_SIG, ROM14_DATA4_SIG,
       ROM14_DATA5_SIG, ROM14_DATA6_SIG, ROM14_DATA7_SIG, ROM14_DATA8_SIG, ROM14_DATA9_SIG,
       ROM14_DATA10_SIG, ROM14_DATA11_SIG, ROM14_DATA12_SIG, ROM14_DATA13_SIG, ROM14_DATA14_SIG,
       ROM14_DATA15_SIG, ROM14_DATA16_SIG, ROM14_DATA17_SIG, ROM14_DATA18_SIG, ROM14_DATA19_SIG,
       ROM14_DATA20_SIG, ROM14_DATA21_SIG, ROM14_DATA22_SIG, ROM14_DATA23_SIG, ROM14_DATA24_SIG, ROM14_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0'); 
signal ROM15_DATA0_SIG, ROM15_DATA1_SIG, ROM15_DATA2_SIG, ROM15_DATA3_SIG, ROM15_DATA4_SIG,
       ROM15_DATA5_SIG, ROM15_DATA6_SIG, ROM15_DATA7_SIG, ROM15_DATA8_SIG, ROM15_DATA9_SIG,
       ROM15_DATA10_SIG, ROM15_DATA11_SIG, ROM15_DATA12_SIG, ROM15_DATA13_SIG, ROM15_DATA14_SIG,
       ROM15_DATA15_SIG, ROM15_DATA16_SIG, ROM15_DATA17_SIG, ROM15_DATA18_SIG, ROM15_DATA19_SIG,
       ROM15_DATA20_SIG, ROM15_DATA21_SIG, ROM15_DATA22_SIG, ROM15_DATA23_SIG, ROM15_DATA24_SIG, ROM15_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0'); 
signal ROM16_DATA0_SIG, ROM16_DATA1_SIG, ROM16_DATA2_SIG, ROM16_DATA3_SIG, ROM16_DATA4_SIG,
       ROM16_DATA5_SIG, ROM16_DATA6_SIG, ROM16_DATA7_SIG, ROM16_DATA8_SIG, ROM16_DATA9_SIG,
       ROM16_DATA10_SIG, ROM16_DATA11_SIG, ROM16_DATA12_SIG, ROM16_DATA13_SIG, ROM16_DATA14_SIG,
       ROM16_DATA15_SIG, ROM16_DATA16_SIG, ROM16_DATA17_SIG, ROM16_DATA18_SIG, ROM16_DATA19_SIG,
       ROM16_DATA20_SIG, ROM16_DATA21_SIG, ROM16_DATA22_SIG, ROM16_DATA23_SIG, ROM16_DATA24_SIG, ROM16_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0'); 
signal ROM17_DATA0_SIG, ROM17_DATA1_SIG, ROM17_DATA2_SIG, ROM17_DATA3_SIG, ROM17_DATA4_SIG,
       ROM17_DATA5_SIG, ROM17_DATA6_SIG, ROM17_DATA7_SIG, ROM17_DATA8_SIG, ROM17_DATA9_SIG,
       ROM17_DATA10_SIG, ROM17_DATA11_SIG, ROM17_DATA12_SIG, ROM17_DATA13_SIG, ROM17_DATA14_SIG,
       ROM17_DATA15_SIG, ROM17_DATA16_SIG, ROM17_DATA17_SIG, ROM17_DATA18_SIG, ROM17_DATA19_SIG,
       ROM17_DATA20_SIG, ROM17_DATA21_SIG, ROM17_DATA22_SIG, ROM17_DATA23_SIG, ROM17_DATA24_SIG, ROM17_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0'); 
signal ROM18_DATA0_SIG, ROM18_DATA1_SIG, ROM18_DATA2_SIG, ROM18_DATA3_SIG, ROM18_DATA4_SIG,
       ROM18_DATA5_SIG, ROM18_DATA6_SIG, ROM18_DATA7_SIG, ROM18_DATA8_SIG, ROM18_DATA9_SIG,
       ROM18_DATA10_SIG, ROM18_DATA11_SIG, ROM18_DATA12_SIG, ROM18_DATA13_SIG, ROM18_DATA14_SIG,
       ROM18_DATA15_SIG, ROM18_DATA16_SIG, ROM18_DATA17_SIG, ROM18_DATA18_SIG, ROM18_DATA19_SIG,
       ROM18_DATA20_SIG, ROM18_DATA21_SIG, ROM18_DATA22_SIG, ROM18_DATA23_SIG, ROM18_DATA24_SIG, ROM18_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0'); 
signal ROM19_DATA0_SIG, ROM19_DATA1_SIG, ROM19_DATA2_SIG, ROM19_DATA3_SIG, ROM19_DATA4_SIG,
       ROM19_DATA5_SIG, ROM19_DATA6_SIG, ROM19_DATA7_SIG, ROM19_DATA8_SIG, ROM19_DATA9_SIG,
       ROM19_DATA10_SIG, ROM19_DATA11_SIG, ROM19_DATA12_SIG, ROM19_DATA13_SIG, ROM19_DATA14_SIG,
       ROM19_DATA15_SIG, ROM19_DATA16_SIG, ROM19_DATA17_SIG, ROM19_DATA18_SIG, ROM19_DATA19_SIG,
       ROM19_DATA20_SIG, ROM19_DATA21_SIG, ROM19_DATA22_SIG, ROM19_DATA23_SIG, ROM19_DATA24_SIG, ROM19_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0'); 
signal ROM20_DATA0_SIG, ROM20_DATA1_SIG, ROM20_DATA2_SIG, ROM20_DATA3_SIG, ROM20_DATA4_SIG,
       ROM20_DATA5_SIG, ROM20_DATA6_SIG, ROM20_DATA7_SIG, ROM20_DATA8_SIG, ROM20_DATA9_SIG,
       ROM20_DATA10_SIG, ROM20_DATA11_SIG, ROM20_DATA12_SIG, ROM20_DATA13_SIG, ROM20_DATA14_SIG,
       ROM20_DATA15_SIG, ROM20_DATA16_SIG, ROM20_DATA17_SIG, ROM20_DATA18_SIG, ROM20_DATA19_SIG,
       ROM20_DATA20_SIG, ROM20_DATA21_SIG, ROM20_DATA22_SIG, ROM20_DATA23_SIG, ROM20_DATA24_SIG, ROM20_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM21_DATA0_SIG, ROM21_DATA1_SIG, ROM21_DATA2_SIG, ROM21_DATA3_SIG, ROM21_DATA4_SIG,
       ROM21_DATA5_SIG, ROM21_DATA6_SIG, ROM21_DATA7_SIG, ROM21_DATA8_SIG, ROM21_DATA9_SIG,
       ROM21_DATA10_SIG, ROM21_DATA11_SIG, ROM21_DATA12_SIG, ROM21_DATA13_SIG, ROM21_DATA14_SIG,
       ROM21_DATA15_SIG, ROM21_DATA16_SIG, ROM21_DATA17_SIG, ROM21_DATA18_SIG, ROM21_DATA19_SIG,
       ROM21_DATA20_SIG, ROM21_DATA21_SIG, ROM21_DATA22_SIG, ROM21_DATA23_SIG, ROM21_DATA24_SIG, ROM21_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM22_DATA0_SIG, ROM22_DATA1_SIG, ROM22_DATA2_SIG, ROM22_DATA3_SIG, ROM22_DATA4_SIG,
       ROM22_DATA5_SIG, ROM22_DATA6_SIG, ROM22_DATA7_SIG, ROM22_DATA8_SIG, ROM22_DATA9_SIG,
       ROM22_DATA10_SIG, ROM22_DATA11_SIG, ROM22_DATA12_SIG, ROM22_DATA13_SIG, ROM22_DATA14_SIG,
       ROM22_DATA15_SIG, ROM22_DATA16_SIG, ROM22_DATA17_SIG, ROM22_DATA18_SIG, ROM22_DATA19_SIG,
       ROM22_DATA20_SIG, ROM22_DATA21_SIG, ROM22_DATA22_SIG, ROM22_DATA23_SIG, ROM22_DATA24_SIG, ROM22_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM23_DATA0_SIG, ROM23_DATA1_SIG, ROM23_DATA2_SIG, ROM23_DATA3_SIG, ROM23_DATA4_SIG,
       ROM23_DATA5_SIG, ROM23_DATA6_SIG, ROM23_DATA7_SIG, ROM23_DATA8_SIG, ROM23_DATA9_SIG,
       ROM23_DATA10_SIG, ROM23_DATA11_SIG, ROM23_DATA12_SIG, ROM23_DATA13_SIG, ROM23_DATA14_SIG,
       ROM23_DATA15_SIG, ROM23_DATA16_SIG, ROM23_DATA17_SIG, ROM23_DATA18_SIG, ROM23_DATA19_SIG,
       ROM23_DATA20_SIG, ROM23_DATA21_SIG, ROM23_DATA22_SIG, ROM23_DATA23_SIG, ROM23_DATA24_SIG, ROM23_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM24_DATA0_SIG, ROM24_DATA1_SIG, ROM24_DATA2_SIG, ROM24_DATA3_SIG, ROM24_DATA4_SIG,
       ROM24_DATA5_SIG, ROM24_DATA6_SIG, ROM24_DATA7_SIG, ROM24_DATA8_SIG, ROM24_DATA9_SIG,
       ROM24_DATA10_SIG, ROM24_DATA11_SIG, ROM24_DATA12_SIG, ROM24_DATA13_SIG, ROM24_DATA14_SIG,
       ROM24_DATA15_SIG, ROM24_DATA16_SIG, ROM24_DATA17_SIG, ROM24_DATA18_SIG, ROM24_DATA19_SIG,
       ROM24_DATA20_SIG, ROM24_DATA21_SIG, ROM24_DATA22_SIG, ROM24_DATA23_SIG, ROM24_DATA24_SIG, ROM24_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM25_DATA0_SIG, ROM25_DATA1_SIG, ROM25_DATA2_SIG, ROM25_DATA3_SIG, ROM25_DATA4_SIG,
       ROM25_DATA5_SIG, ROM25_DATA6_SIG, ROM25_DATA7_SIG, ROM25_DATA8_SIG, ROM25_DATA9_SIG,
       ROM25_DATA10_SIG, ROM25_DATA11_SIG, ROM25_DATA12_SIG, ROM25_DATA13_SIG, ROM25_DATA14_SIG,
       ROM25_DATA15_SIG, ROM25_DATA16_SIG, ROM25_DATA17_SIG, ROM25_DATA18_SIG, ROM25_DATA19_SIG,
       ROM25_DATA20_SIG, ROM25_DATA21_SIG, ROM25_DATA22_SIG, ROM25_DATA23_SIG, ROM25_DATA24_SIG, ROM25_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM26_DATA0_SIG, ROM26_DATA1_SIG, ROM26_DATA2_SIG, ROM26_DATA3_SIG, ROM26_DATA4_SIG,
       ROM26_DATA5_SIG, ROM26_DATA6_SIG, ROM26_DATA7_SIG, ROM26_DATA8_SIG, ROM26_DATA9_SIG,
       ROM26_DATA10_SIG, ROM26_DATA11_SIG, ROM26_DATA12_SIG, ROM26_DATA13_SIG, ROM26_DATA14_SIG,
       ROM26_DATA15_SIG, ROM26_DATA16_SIG, ROM26_DATA17_SIG, ROM26_DATA18_SIG, ROM26_DATA19_SIG,
       ROM26_DATA20_SIG, ROM26_DATA21_SIG, ROM26_DATA22_SIG, ROM26_DATA23_SIG, ROM26_DATA24_SIG, ROM26_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM27_DATA0_SIG, ROM27_DATA1_SIG, ROM27_DATA2_SIG, ROM27_DATA3_SIG, ROM27_DATA4_SIG,
       ROM27_DATA5_SIG, ROM27_DATA6_SIG, ROM27_DATA7_SIG, ROM27_DATA8_SIG, ROM27_DATA9_SIG,
       ROM27_DATA10_SIG, ROM27_DATA11_SIG, ROM27_DATA12_SIG, ROM27_DATA13_SIG, ROM27_DATA14_SIG,
       ROM27_DATA15_SIG, ROM27_DATA16_SIG, ROM27_DATA17_SIG, ROM27_DATA18_SIG, ROM27_DATA19_SIG,
       ROM27_DATA20_SIG, ROM27_DATA21_SIG, ROM27_DATA22_SIG, ROM27_DATA23_SIG, ROM27_DATA24_SIG, ROM27_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM28_DATA0_SIG, ROM28_DATA1_SIG, ROM28_DATA2_SIG, ROM28_DATA3_SIG, ROM28_DATA4_SIG,
       ROM28_DATA5_SIG, ROM28_DATA6_SIG, ROM28_DATA7_SIG, ROM28_DATA8_SIG, ROM28_DATA9_SIG,
       ROM28_DATA10_SIG, ROM28_DATA11_SIG, ROM28_DATA12_SIG, ROM28_DATA13_SIG, ROM28_DATA14_SIG,
       ROM28_DATA15_SIG, ROM28_DATA16_SIG, ROM28_DATA17_SIG, ROM28_DATA18_SIG, ROM28_DATA19_SIG,
       ROM28_DATA20_SIG, ROM28_DATA21_SIG, ROM28_DATA22_SIG, ROM28_DATA23_SIG, ROM28_DATA24_SIG, ROM28_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM29_DATA0_SIG, ROM29_DATA1_SIG, ROM29_DATA2_SIG, ROM29_DATA3_SIG, ROM29_DATA4_SIG,
       ROM29_DATA5_SIG, ROM29_DATA6_SIG, ROM29_DATA7_SIG, ROM29_DATA8_SIG, ROM29_DATA9_SIG,
       ROM29_DATA10_SIG, ROM29_DATA11_SIG, ROM29_DATA12_SIG, ROM29_DATA13_SIG, ROM29_DATA14_SIG,
       ROM29_DATA15_SIG, ROM29_DATA16_SIG, ROM29_DATA17_SIG, ROM29_DATA18_SIG, ROM29_DATA19_SIG,
       ROM29_DATA20_SIG, ROM29_DATA21_SIG, ROM29_DATA22_SIG, ROM29_DATA23_SIG, ROM29_DATA24_SIG, ROM29_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM30_DATA0_SIG, ROM30_DATA1_SIG, ROM30_DATA2_SIG, ROM30_DATA3_SIG, ROM30_DATA4_SIG,
       ROM30_DATA5_SIG, ROM30_DATA6_SIG, ROM30_DATA7_SIG, ROM30_DATA8_SIG, ROM30_DATA9_SIG,
       ROM30_DATA10_SIG, ROM30_DATA11_SIG, ROM30_DATA12_SIG, ROM30_DATA13_SIG, ROM30_DATA14_SIG,
       ROM30_DATA15_SIG, ROM30_DATA16_SIG, ROM30_DATA17_SIG, ROM30_DATA18_SIG, ROM30_DATA19_SIG,
       ROM30_DATA20_SIG, ROM30_DATA21_SIG, ROM30_DATA22_SIG, ROM30_DATA23_SIG, ROM30_DATA24_SIG, ROM30_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
signal ROM31_DATA0_SIG, ROM31_DATA1_SIG, ROM31_DATA2_SIG, ROM31_DATA3_SIG, ROM31_DATA4_SIG,
       ROM31_DATA5_SIG, ROM31_DATA6_SIG, ROM31_DATA7_SIG, ROM31_DATA8_SIG, ROM31_DATA9_SIG,
       ROM31_DATA10_SIG, ROM31_DATA11_SIG, ROM31_DATA12_SIG, ROM31_DATA13_SIG, ROM31_DATA14_SIG,
       ROM31_DATA15_SIG, ROM31_DATA16_SIG, ROM31_DATA17_SIG, ROM31_DATA18_SIG, ROM31_DATA19_SIG,
       ROM31_DATA20_SIG, ROM31_DATA21_SIG, ROM31_DATA22_SIG, ROM31_DATA23_SIG, ROM31_DATA24_SIG, ROM31_DATA25_SIG : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
begin

DIN0_SIG <= DIN0;
DIN1_SIG <= DIN1;
DIN2_SIG <= DIN2;
DIN3_SIG <= DIN3;
DIN4_SIG <= DIN4;

DSP_BLOCK0_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM0_DATA0_SIG,
    PE01_COEF => ROM0_DATA1_SIG,
    PE02_COEF => ROM0_DATA2_SIG,
    PE03_COEF => ROM0_DATA3_SIG,
    PE04_COEF => ROM0_DATA4_SIG,
    PE10_COEF => ROM0_DATA5_SIG,
    PE11_COEF => ROM0_DATA6_SIG,
    PE12_COEF => ROM0_DATA7_SIG,
    PE13_COEF => ROM0_DATA8_SIG,
    PE14_COEF => ROM0_DATA9_SIG,
    PE20_COEF => ROM0_DATA10_SIG,
    PE21_COEF => ROM0_DATA11_SIG,
    PE22_COEF => ROM0_DATA12_SIG,
    PE23_COEF => ROM0_DATA13_SIG,
    PE24_COEF => ROM0_DATA14_SIG,
    PE30_COEF => ROM0_DATA15_SIG,
    PE31_COEF => ROM0_DATA16_SIG,
    PE32_COEF => ROM0_DATA17_SIG,
    PE33_COEF => ROM0_DATA18_SIG,
    PE34_COEF => ROM0_DATA19_SIG,
    PE40_COEF => ROM0_DATA20_SIG,
    PE41_COEF => ROM0_DATA21_SIG,
    PE42_COEF => ROM0_DATA22_SIG,
    PE43_COEF => ROM0_DATA23_SIG,
    PE44_COEF => ROM0_DATA24_SIG,
    BIAS      => ROM0_DATA25_SIG,
    DOUT      => DOUT0_SIG
);

DSP_BLOCK1_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM1_DATA0_SIG,
    PE01_COEF => ROM1_DATA1_SIG,
    PE02_COEF => ROM1_DATA2_SIG,
    PE03_COEF => ROM1_DATA3_SIG,
    PE04_COEF => ROM1_DATA4_SIG,
    PE10_COEF => ROM1_DATA5_SIG,
    PE11_COEF => ROM1_DATA6_SIG,
    PE12_COEF => ROM1_DATA7_SIG,
    PE13_COEF => ROM1_DATA8_SIG,
    PE14_COEF => ROM1_DATA9_SIG,
    PE20_COEF => ROM1_DATA10_SIG,
    PE21_COEF => ROM1_DATA11_SIG,
    PE22_COEF => ROM1_DATA12_SIG,
    PE23_COEF => ROM1_DATA13_SIG,
    PE24_COEF => ROM1_DATA14_SIG,
    PE30_COEF => ROM1_DATA15_SIG,
    PE31_COEF => ROM1_DATA16_SIG,
    PE32_COEF => ROM1_DATA17_SIG,
    PE33_COEF => ROM1_DATA18_SIG,
    PE34_COEF => ROM1_DATA19_SIG,
    PE40_COEF => ROM1_DATA20_SIG,
    PE41_COEF => ROM1_DATA21_SIG,
    PE42_COEF => ROM1_DATA22_SIG,
    PE43_COEF => ROM1_DATA23_SIG,
    PE44_COEF => ROM1_DATA24_SIG,
    BIAS      => ROM1_DATA25_SIG,
    DOUT      => DOUT1_SIG
);

DSP_BLOCK2_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM2_DATA0_SIG,
    PE01_COEF => ROM2_DATA1_SIG,
    PE02_COEF => ROM2_DATA2_SIG,
    PE03_COEF => ROM2_DATA3_SIG,
    PE04_COEF => ROM2_DATA4_SIG,
    PE10_COEF => ROM2_DATA5_SIG,
    PE11_COEF => ROM2_DATA6_SIG,
    PE12_COEF => ROM2_DATA7_SIG,
    PE13_COEF => ROM2_DATA8_SIG,
    PE14_COEF => ROM2_DATA9_SIG,
    PE20_COEF => ROM2_DATA10_SIG,
    PE21_COEF => ROM2_DATA11_SIG,
    PE22_COEF => ROM2_DATA12_SIG,
    PE23_COEF => ROM2_DATA13_SIG,
    PE24_COEF => ROM2_DATA14_SIG,
    PE30_COEF => ROM2_DATA15_SIG,
    PE31_COEF => ROM2_DATA16_SIG,
    PE32_COEF => ROM2_DATA17_SIG,
    PE33_COEF => ROM2_DATA18_SIG,
    PE34_COEF => ROM2_DATA19_SIG,
    PE40_COEF => ROM2_DATA20_SIG,
    PE41_COEF => ROM2_DATA21_SIG,
    PE42_COEF => ROM2_DATA22_SIG,
    PE43_COEF => ROM2_DATA23_SIG,
    PE44_COEF => ROM2_DATA24_SIG,
    BIAS      => ROM2_DATA25_SIG,
    DOUT      => DOUT2_SIG
);

DSP_BLOCK3_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM3_DATA0_SIG,
    PE01_COEF => ROM3_DATA1_SIG,
    PE02_COEF => ROM3_DATA2_SIG,
    PE03_COEF => ROM3_DATA3_SIG,
    PE04_COEF => ROM3_DATA4_SIG,
    PE10_COEF => ROM3_DATA5_SIG,
    PE11_COEF => ROM3_DATA6_SIG,
    PE12_COEF => ROM3_DATA7_SIG,
    PE13_COEF => ROM3_DATA8_SIG,
    PE14_COEF => ROM3_DATA9_SIG,
    PE20_COEF => ROM3_DATA10_SIG,
    PE21_COEF => ROM3_DATA11_SIG,
    PE22_COEF => ROM3_DATA12_SIG,
    PE23_COEF => ROM3_DATA13_SIG,
    PE24_COEF => ROM3_DATA14_SIG,
    PE30_COEF => ROM3_DATA15_SIG,
    PE31_COEF => ROM3_DATA16_SIG,
    PE32_COEF => ROM3_DATA17_SIG,
    PE33_COEF => ROM3_DATA18_SIG,
    PE34_COEF => ROM3_DATA19_SIG,
    PE40_COEF => ROM3_DATA20_SIG,
    PE41_COEF => ROM3_DATA21_SIG,
    PE42_COEF => ROM3_DATA22_SIG,
    PE43_COEF => ROM3_DATA23_SIG,
    PE44_COEF => ROM3_DATA24_SIG,
    BIAS      => ROM3_DATA25_SIG,
    DOUT      => DOUT3_SIG
);

DSP_BLOCK4_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM4_DATA0_SIG,
    PE01_COEF => ROM4_DATA1_SIG,
    PE02_COEF => ROM4_DATA2_SIG,
    PE03_COEF => ROM4_DATA3_SIG,
    PE04_COEF => ROM4_DATA4_SIG,
    PE10_COEF => ROM4_DATA5_SIG,
    PE11_COEF => ROM4_DATA6_SIG,
    PE12_COEF => ROM4_DATA7_SIG,
    PE13_COEF => ROM4_DATA8_SIG,
    PE14_COEF => ROM4_DATA9_SIG,
    PE20_COEF => ROM4_DATA10_SIG,
    PE21_COEF => ROM4_DATA11_SIG,
    PE22_COEF => ROM4_DATA12_SIG,
    PE23_COEF => ROM4_DATA13_SIG,
    PE24_COEF => ROM4_DATA14_SIG,
    PE30_COEF => ROM4_DATA15_SIG,
    PE31_COEF => ROM4_DATA16_SIG,
    PE32_COEF => ROM4_DATA17_SIG,
    PE33_COEF => ROM4_DATA18_SIG,
    PE34_COEF => ROM4_DATA19_SIG,
    PE40_COEF => ROM4_DATA20_SIG,
    PE41_COEF => ROM4_DATA21_SIG,
    PE42_COEF => ROM4_DATA22_SIG,
    PE43_COEF => ROM4_DATA23_SIG,
    PE44_COEF => ROM4_DATA24_SIG,
    BIAS      => ROM4_DATA25_SIG,
    DOUT      => DOUT4_SIG
);

DSP_BLOCK5_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM5_DATA0_SIG,
    PE01_COEF => ROM5_DATA1_SIG,
    PE02_COEF => ROM5_DATA2_SIG,
    PE03_COEF => ROM5_DATA3_SIG,
    PE04_COEF => ROM5_DATA4_SIG,
    PE10_COEF => ROM5_DATA5_SIG,
    PE11_COEF => ROM5_DATA6_SIG,
    PE12_COEF => ROM5_DATA7_SIG,
    PE13_COEF => ROM5_DATA8_SIG,
    PE14_COEF => ROM5_DATA9_SIG,
    PE20_COEF => ROM5_DATA10_SIG,
    PE21_COEF => ROM5_DATA11_SIG,
    PE22_COEF => ROM5_DATA12_SIG,
    PE23_COEF => ROM5_DATA13_SIG,
    PE24_COEF => ROM5_DATA14_SIG,
    PE30_COEF => ROM5_DATA15_SIG,
    PE31_COEF => ROM5_DATA16_SIG,
    PE32_COEF => ROM5_DATA17_SIG,
    PE33_COEF => ROM5_DATA18_SIG,
    PE34_COEF => ROM5_DATA19_SIG,
    PE40_COEF => ROM5_DATA20_SIG,
    PE41_COEF => ROM5_DATA21_SIG,
    PE42_COEF => ROM5_DATA22_SIG,
    PE43_COEF => ROM5_DATA23_SIG,
    PE44_COEF => ROM5_DATA24_SIG,
    BIAS      => ROM5_DATA25_SIG,
    DOUT      => DOUT5_SIG
);

DSP_BLOCK6_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM6_DATA0_SIG,
    PE01_COEF => ROM6_DATA1_SIG,
    PE02_COEF => ROM6_DATA2_SIG,
    PE03_COEF => ROM6_DATA3_SIG,
    PE04_COEF => ROM6_DATA4_SIG,
    PE10_COEF => ROM6_DATA5_SIG,
    PE11_COEF => ROM6_DATA6_SIG,
    PE12_COEF => ROM6_DATA7_SIG,
    PE13_COEF => ROM6_DATA8_SIG,
    PE14_COEF => ROM6_DATA9_SIG,
    PE20_COEF => ROM6_DATA10_SIG,
    PE21_COEF => ROM6_DATA11_SIG,
    PE22_COEF => ROM6_DATA12_SIG,
    PE23_COEF => ROM6_DATA13_SIG,
    PE24_COEF => ROM6_DATA14_SIG,
    PE30_COEF => ROM6_DATA15_SIG,
    PE31_COEF => ROM6_DATA16_SIG,
    PE32_COEF => ROM6_DATA17_SIG,
    PE33_COEF => ROM6_DATA18_SIG,
    PE34_COEF => ROM6_DATA19_SIG,
    PE40_COEF => ROM6_DATA20_SIG,
    PE41_COEF => ROM6_DATA21_SIG,
    PE42_COEF => ROM6_DATA22_SIG,
    PE43_COEF => ROM6_DATA23_SIG,
    PE44_COEF => ROM6_DATA24_SIG,
    BIAS      => ROM6_DATA25_SIG,
    DOUT      => DOUT6_SIG
);

DSP_BLOCK7_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM7_DATA0_SIG,
    PE01_COEF => ROM7_DATA1_SIG,
    PE02_COEF => ROM7_DATA2_SIG,
    PE03_COEF => ROM7_DATA3_SIG,
    PE04_COEF => ROM7_DATA4_SIG,
    PE10_COEF => ROM7_DATA5_SIG,
    PE11_COEF => ROM7_DATA6_SIG,
    PE12_COEF => ROM7_DATA7_SIG,
    PE13_COEF => ROM7_DATA8_SIG,
    PE14_COEF => ROM7_DATA9_SIG,
    PE20_COEF => ROM7_DATA10_SIG,
    PE21_COEF => ROM7_DATA11_SIG,
    PE22_COEF => ROM7_DATA12_SIG,
    PE23_COEF => ROM7_DATA13_SIG,
    PE24_COEF => ROM7_DATA14_SIG,
    PE30_COEF => ROM7_DATA15_SIG,
    PE31_COEF => ROM7_DATA16_SIG,
    PE32_COEF => ROM7_DATA17_SIG,
    PE33_COEF => ROM7_DATA18_SIG,
    PE34_COEF => ROM7_DATA19_SIG,
    PE40_COEF => ROM7_DATA20_SIG,
    PE41_COEF => ROM7_DATA21_SIG,
    PE42_COEF => ROM7_DATA22_SIG,
    PE43_COEF => ROM7_DATA23_SIG,
    PE44_COEF => ROM7_DATA24_SIG,
    BIAS      => ROM7_DATA25_SIG,
    DOUT      => DOUT7_SIG
);

DSP_BLOCK8_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM8_DATA0_SIG,
    PE01_COEF => ROM8_DATA1_SIG,
    PE02_COEF => ROM8_DATA2_SIG,
    PE03_COEF => ROM8_DATA3_SIG,
    PE04_COEF => ROM8_DATA4_SIG,
    PE10_COEF => ROM8_DATA5_SIG,
    PE11_COEF => ROM8_DATA6_SIG,
    PE12_COEF => ROM8_DATA7_SIG,
    PE13_COEF => ROM8_DATA8_SIG,
    PE14_COEF => ROM8_DATA9_SIG,
    PE20_COEF => ROM8_DATA10_SIG,
    PE21_COEF => ROM8_DATA11_SIG,
    PE22_COEF => ROM8_DATA12_SIG,
    PE23_COEF => ROM8_DATA13_SIG,
    PE24_COEF => ROM8_DATA14_SIG,
    PE30_COEF => ROM8_DATA15_SIG,
    PE31_COEF => ROM8_DATA16_SIG,
    PE32_COEF => ROM8_DATA17_SIG,
    PE33_COEF => ROM8_DATA18_SIG,
    PE34_COEF => ROM8_DATA19_SIG,
    PE40_COEF => ROM8_DATA20_SIG,
    PE41_COEF => ROM8_DATA21_SIG,
    PE42_COEF => ROM8_DATA22_SIG,
    PE43_COEF => ROM8_DATA23_SIG,
    PE44_COEF => ROM8_DATA24_SIG,
    BIAS      => ROM8_DATA25_SIG,
    DOUT      => DOUT8_SIG
);

DSP_BLOCK9_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM9_DATA0_SIG,
    PE01_COEF => ROM9_DATA1_SIG,
    PE02_COEF => ROM9_DATA2_SIG,
    PE03_COEF => ROM9_DATA3_SIG,
    PE04_COEF => ROM9_DATA4_SIG,
    PE10_COEF => ROM9_DATA5_SIG,
    PE11_COEF => ROM9_DATA6_SIG,
    PE12_COEF => ROM9_DATA7_SIG,
    PE13_COEF => ROM9_DATA8_SIG,
    PE14_COEF => ROM9_DATA9_SIG,
    PE20_COEF => ROM9_DATA10_SIG,
    PE21_COEF => ROM9_DATA11_SIG,
    PE22_COEF => ROM9_DATA12_SIG,
    PE23_COEF => ROM9_DATA13_SIG,
    PE24_COEF => ROM9_DATA14_SIG,
    PE30_COEF => ROM9_DATA15_SIG,
    PE31_COEF => ROM9_DATA16_SIG,
    PE32_COEF => ROM9_DATA17_SIG,
    PE33_COEF => ROM9_DATA18_SIG,
    PE34_COEF => ROM9_DATA19_SIG,
    PE40_COEF => ROM9_DATA20_SIG,
    PE41_COEF => ROM9_DATA21_SIG,
    PE42_COEF => ROM9_DATA22_SIG,
    PE43_COEF => ROM9_DATA23_SIG,
    PE44_COEF => ROM9_DATA24_SIG,
    BIAS      => ROM9_DATA25_SIG,
    DOUT      => DOUT9_SIG
);

DSP_BLOCK10_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM10_DATA0_SIG,
    PE01_COEF => ROM10_DATA1_SIG,
    PE02_COEF => ROM10_DATA2_SIG,
    PE03_COEF => ROM10_DATA3_SIG,
    PE04_COEF => ROM10_DATA4_SIG,
    PE10_COEF => ROM10_DATA5_SIG,
    PE11_COEF => ROM10_DATA6_SIG,
    PE12_COEF => ROM10_DATA7_SIG,
    PE13_COEF => ROM10_DATA8_SIG,
    PE14_COEF => ROM10_DATA9_SIG,
    PE20_COEF => ROM10_DATA10_SIG,
    PE21_COEF => ROM10_DATA11_SIG,
    PE22_COEF => ROM10_DATA12_SIG,
    PE23_COEF => ROM10_DATA13_SIG,
    PE24_COEF => ROM10_DATA14_SIG,
    PE30_COEF => ROM10_DATA15_SIG,
    PE31_COEF => ROM10_DATA16_SIG,
    PE32_COEF => ROM10_DATA17_SIG,
    PE33_COEF => ROM10_DATA18_SIG,
    PE34_COEF => ROM10_DATA19_SIG,
    PE40_COEF => ROM10_DATA20_SIG,
    PE41_COEF => ROM10_DATA21_SIG,
    PE42_COEF => ROM10_DATA22_SIG,
    PE43_COEF => ROM10_DATA23_SIG,
    PE44_COEF => ROM10_DATA24_SIG,
    BIAS      => ROM10_DATA25_SIG,
    DOUT      => DOUT10_SIG
);

DSP_BLOCK11_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM11_DATA0_SIG,
    PE01_COEF => ROM11_DATA1_SIG,
    PE02_COEF => ROM11_DATA2_SIG,
    PE03_COEF => ROM11_DATA3_SIG,
    PE04_COEF => ROM11_DATA4_SIG,
    PE10_COEF => ROM11_DATA5_SIG,
    PE11_COEF => ROM11_DATA6_SIG,
    PE12_COEF => ROM11_DATA7_SIG,
    PE13_COEF => ROM11_DATA8_SIG,
    PE14_COEF => ROM11_DATA9_SIG,
    PE20_COEF => ROM11_DATA10_SIG,
    PE21_COEF => ROM11_DATA11_SIG,
    PE22_COEF => ROM11_DATA12_SIG,
    PE23_COEF => ROM11_DATA13_SIG,
    PE24_COEF => ROM11_DATA14_SIG,
    PE30_COEF => ROM11_DATA15_SIG,
    PE31_COEF => ROM11_DATA16_SIG,
    PE32_COEF => ROM11_DATA17_SIG,
    PE33_COEF => ROM11_DATA18_SIG,
    PE34_COEF => ROM11_DATA19_SIG,
    PE40_COEF => ROM11_DATA20_SIG,
    PE41_COEF => ROM11_DATA21_SIG,
    PE42_COEF => ROM11_DATA22_SIG,
    PE43_COEF => ROM11_DATA23_SIG,
    PE44_COEF => ROM11_DATA24_SIG,
    BIAS      => ROM11_DATA25_SIG,
    DOUT      => DOUT11_SIG
);

DSP_BLOCK12_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM12_DATA0_SIG,
    PE01_COEF => ROM12_DATA1_SIG,
    PE02_COEF => ROM12_DATA2_SIG,
    PE03_COEF => ROM12_DATA3_SIG,
    PE04_COEF => ROM12_DATA4_SIG,
    PE10_COEF => ROM12_DATA5_SIG,
    PE11_COEF => ROM12_DATA6_SIG,
    PE12_COEF => ROM12_DATA7_SIG,
    PE13_COEF => ROM12_DATA8_SIG,
    PE14_COEF => ROM12_DATA9_SIG,
    PE20_COEF => ROM12_DATA10_SIG,
    PE21_COEF => ROM12_DATA11_SIG,
    PE22_COEF => ROM12_DATA12_SIG,
    PE23_COEF => ROM12_DATA13_SIG,
    PE24_COEF => ROM12_DATA14_SIG,
    PE30_COEF => ROM12_DATA15_SIG,
    PE31_COEF => ROM12_DATA16_SIG,
    PE32_COEF => ROM12_DATA17_SIG,
    PE33_COEF => ROM12_DATA18_SIG,
    PE34_COEF => ROM12_DATA19_SIG,
    PE40_COEF => ROM12_DATA20_SIG,
    PE41_COEF => ROM12_DATA21_SIG,
    PE42_COEF => ROM12_DATA22_SIG,
    PE43_COEF => ROM12_DATA23_SIG,
    PE44_COEF => ROM12_DATA24_SIG,
    BIAS      => ROM12_DATA25_SIG,
    DOUT      => DOUT12_SIG
);

DSP_BLOCK13_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM13_DATA0_SIG,
    PE01_COEF => ROM13_DATA1_SIG,
    PE02_COEF => ROM13_DATA2_SIG,
    PE03_COEF => ROM13_DATA3_SIG,
    PE04_COEF => ROM13_DATA4_SIG,
    PE10_COEF => ROM13_DATA5_SIG,
    PE11_COEF => ROM13_DATA6_SIG,
    PE12_COEF => ROM13_DATA7_SIG,
    PE13_COEF => ROM13_DATA8_SIG,
    PE14_COEF => ROM13_DATA9_SIG,
    PE20_COEF => ROM13_DATA10_SIG,
    PE21_COEF => ROM13_DATA11_SIG,
    PE22_COEF => ROM13_DATA12_SIG,
    PE23_COEF => ROM13_DATA13_SIG,
    PE24_COEF => ROM13_DATA14_SIG,
    PE30_COEF => ROM13_DATA15_SIG,
    PE31_COEF => ROM13_DATA16_SIG,
    PE32_COEF => ROM13_DATA17_SIG,
    PE33_COEF => ROM13_DATA18_SIG,
    PE34_COEF => ROM13_DATA19_SIG,
    PE40_COEF => ROM13_DATA20_SIG,
    PE41_COEF => ROM13_DATA21_SIG,
    PE42_COEF => ROM13_DATA22_SIG,
    PE43_COEF => ROM13_DATA23_SIG,
    PE44_COEF => ROM13_DATA24_SIG,
    BIAS      => ROM13_DATA25_SIG,
    DOUT      => DOUT13_SIG
);

DSP_BLOCK14_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM14_DATA0_SIG,
    PE01_COEF => ROM14_DATA1_SIG,
    PE02_COEF => ROM14_DATA2_SIG,
    PE03_COEF => ROM14_DATA3_SIG,
    PE04_COEF => ROM14_DATA4_SIG,
    PE10_COEF => ROM14_DATA5_SIG,
    PE11_COEF => ROM14_DATA6_SIG,
    PE12_COEF => ROM14_DATA7_SIG,
    PE13_COEF => ROM14_DATA8_SIG,
    PE14_COEF => ROM14_DATA9_SIG,
    PE20_COEF => ROM14_DATA10_SIG,
    PE21_COEF => ROM14_DATA11_SIG,
    PE22_COEF => ROM14_DATA12_SIG,
    PE23_COEF => ROM14_DATA13_SIG,
    PE24_COEF => ROM14_DATA14_SIG,
    PE30_COEF => ROM14_DATA15_SIG,
    PE31_COEF => ROM14_DATA16_SIG,
    PE32_COEF => ROM14_DATA17_SIG,
    PE33_COEF => ROM14_DATA18_SIG,
    PE34_COEF => ROM14_DATA19_SIG,
    PE40_COEF => ROM14_DATA20_SIG,
    PE41_COEF => ROM14_DATA21_SIG,
    PE42_COEF => ROM14_DATA22_SIG,
    PE43_COEF => ROM14_DATA23_SIG,
    PE44_COEF => ROM14_DATA24_SIG,
    BIAS      => ROM14_DATA25_SIG,
    DOUT      => DOUT14_SIG
);

DSP_BLOCK15_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM15_DATA0_SIG,
    PE01_COEF => ROM15_DATA1_SIG,
    PE02_COEF => ROM15_DATA2_SIG,
    PE03_COEF => ROM15_DATA3_SIG,
    PE04_COEF => ROM15_DATA4_SIG,
    PE10_COEF => ROM15_DATA5_SIG,
    PE11_COEF => ROM15_DATA6_SIG,
    PE12_COEF => ROM15_DATA7_SIG,
    PE13_COEF => ROM15_DATA8_SIG,
    PE14_COEF => ROM15_DATA9_SIG,
    PE20_COEF => ROM15_DATA10_SIG,
    PE21_COEF => ROM15_DATA11_SIG,
    PE22_COEF => ROM15_DATA12_SIG,
    PE23_COEF => ROM15_DATA13_SIG,
    PE24_COEF => ROM15_DATA14_SIG,
    PE30_COEF => ROM15_DATA15_SIG,
    PE31_COEF => ROM15_DATA16_SIG,
    PE32_COEF => ROM15_DATA17_SIG,
    PE33_COEF => ROM15_DATA18_SIG,
    PE34_COEF => ROM15_DATA19_SIG,
    PE40_COEF => ROM15_DATA20_SIG,
    PE41_COEF => ROM15_DATA21_SIG,
    PE42_COEF => ROM15_DATA22_SIG,
    PE43_COEF => ROM15_DATA23_SIG,
    PE44_COEF => ROM15_DATA24_SIG,
    BIAS      => ROM15_DATA25_SIG,
    DOUT      => DOUT15_SIG
);

DSP_BLOCK16_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM16_DATA0_SIG,
    PE01_COEF => ROM16_DATA1_SIG,
    PE02_COEF => ROM16_DATA2_SIG,
    PE03_COEF => ROM16_DATA3_SIG,
    PE04_COEF => ROM16_DATA4_SIG,
    PE10_COEF => ROM16_DATA5_SIG,
    PE11_COEF => ROM16_DATA6_SIG,
    PE12_COEF => ROM16_DATA7_SIG,
    PE13_COEF => ROM16_DATA8_SIG,
    PE14_COEF => ROM16_DATA9_SIG,
    PE20_COEF => ROM16_DATA10_SIG,
    PE21_COEF => ROM16_DATA11_SIG,
    PE22_COEF => ROM16_DATA12_SIG,
    PE23_COEF => ROM16_DATA13_SIG,
    PE24_COEF => ROM16_DATA14_SIG,
    PE30_COEF => ROM16_DATA15_SIG,
    PE31_COEF => ROM16_DATA16_SIG,
    PE32_COEF => ROM16_DATA17_SIG,
    PE33_COEF => ROM16_DATA18_SIG,
    PE34_COEF => ROM16_DATA19_SIG,
    PE40_COEF => ROM16_DATA20_SIG,
    PE41_COEF => ROM16_DATA21_SIG,
    PE42_COEF => ROM16_DATA22_SIG,
    PE43_COEF => ROM16_DATA23_SIG,
    PE44_COEF => ROM16_DATA24_SIG,
    BIAS      => ROM16_DATA25_SIG,
    DOUT      => DOUT16_SIG
);

DSP_BLOCK17_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM17_DATA0_SIG,
    PE01_COEF => ROM17_DATA1_SIG,
    PE02_COEF => ROM17_DATA2_SIG,
    PE03_COEF => ROM17_DATA3_SIG,
    PE04_COEF => ROM17_DATA4_SIG,
    PE10_COEF => ROM17_DATA5_SIG,
    PE11_COEF => ROM17_DATA6_SIG,
    PE12_COEF => ROM17_DATA7_SIG,
    PE13_COEF => ROM17_DATA8_SIG,
    PE14_COEF => ROM17_DATA9_SIG,
    PE20_COEF => ROM17_DATA10_SIG,
    PE21_COEF => ROM17_DATA11_SIG,
    PE22_COEF => ROM17_DATA12_SIG,
    PE23_COEF => ROM17_DATA13_SIG,
    PE24_COEF => ROM17_DATA14_SIG,
    PE30_COEF => ROM17_DATA15_SIG,
    PE31_COEF => ROM17_DATA16_SIG,
    PE32_COEF => ROM17_DATA17_SIG,
    PE33_COEF => ROM17_DATA18_SIG,
    PE34_COEF => ROM17_DATA19_SIG,
    PE40_COEF => ROM17_DATA20_SIG,
    PE41_COEF => ROM17_DATA21_SIG,
    PE42_COEF => ROM17_DATA22_SIG,
    PE43_COEF => ROM17_DATA23_SIG,
    PE44_COEF => ROM17_DATA24_SIG,
    BIAS      => ROM17_DATA25_SIG,
    DOUT      => DOUT17_SIG
);

DSP_BLOCK18_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM18_DATA0_SIG,
    PE01_COEF => ROM18_DATA1_SIG,
    PE02_COEF => ROM18_DATA2_SIG,
    PE03_COEF => ROM18_DATA3_SIG,
    PE04_COEF => ROM18_DATA4_SIG,
    PE10_COEF => ROM18_DATA5_SIG,
    PE11_COEF => ROM18_DATA6_SIG,
    PE12_COEF => ROM18_DATA7_SIG,
    PE13_COEF => ROM18_DATA8_SIG,
    PE14_COEF => ROM18_DATA9_SIG,
    PE20_COEF => ROM18_DATA10_SIG,
    PE21_COEF => ROM18_DATA11_SIG,
    PE22_COEF => ROM18_DATA12_SIG,
    PE23_COEF => ROM18_DATA13_SIG,
    PE24_COEF => ROM18_DATA14_SIG,
    PE30_COEF => ROM18_DATA15_SIG,
    PE31_COEF => ROM18_DATA16_SIG,
    PE32_COEF => ROM18_DATA17_SIG,
    PE33_COEF => ROM18_DATA18_SIG,
    PE34_COEF => ROM18_DATA19_SIG,
    PE40_COEF => ROM18_DATA20_SIG,
    PE41_COEF => ROM18_DATA21_SIG,
    PE42_COEF => ROM18_DATA22_SIG,
    PE43_COEF => ROM18_DATA23_SIG,
    PE44_COEF => ROM18_DATA24_SIG,
    BIAS      => ROM18_DATA25_SIG,
    DOUT      => DOUT18_SIG
);

DSP_BLOCK19_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM19_DATA0_SIG,
    PE01_COEF => ROM19_DATA1_SIG,
    PE02_COEF => ROM19_DATA2_SIG,
    PE03_COEF => ROM19_DATA3_SIG,
    PE04_COEF => ROM19_DATA4_SIG,
    PE10_COEF => ROM19_DATA5_SIG,
    PE11_COEF => ROM19_DATA6_SIG,
    PE12_COEF => ROM19_DATA7_SIG,
    PE13_COEF => ROM19_DATA8_SIG,
    PE14_COEF => ROM19_DATA9_SIG,
    PE20_COEF => ROM19_DATA10_SIG,
    PE21_COEF => ROM19_DATA11_SIG,
    PE22_COEF => ROM19_DATA12_SIG,
    PE23_COEF => ROM19_DATA13_SIG,
    PE24_COEF => ROM19_DATA14_SIG,
    PE30_COEF => ROM19_DATA15_SIG,
    PE31_COEF => ROM19_DATA16_SIG,
    PE32_COEF => ROM19_DATA17_SIG,
    PE33_COEF => ROM19_DATA18_SIG,
    PE34_COEF => ROM19_DATA19_SIG,
    PE40_COEF => ROM19_DATA20_SIG,
    PE41_COEF => ROM19_DATA21_SIG,
    PE42_COEF => ROM19_DATA22_SIG,
    PE43_COEF => ROM19_DATA23_SIG,
    PE44_COEF => ROM19_DATA24_SIG,
    BIAS      => ROM19_DATA25_SIG,
    DOUT      => DOUT19_SIG
);

DSP_BLOCK20_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM20_DATA0_SIG,
    PE01_COEF => ROM20_DATA1_SIG,
    PE02_COEF => ROM20_DATA2_SIG,
    PE03_COEF => ROM20_DATA3_SIG,
    PE04_COEF => ROM20_DATA4_SIG,
    PE10_COEF => ROM20_DATA5_SIG,
    PE11_COEF => ROM20_DATA6_SIG,
    PE12_COEF => ROM20_DATA7_SIG,
    PE13_COEF => ROM20_DATA8_SIG,
    PE14_COEF => ROM20_DATA9_SIG,
    PE20_COEF => ROM20_DATA10_SIG,
    PE21_COEF => ROM20_DATA11_SIG,
    PE22_COEF => ROM20_DATA12_SIG,
    PE23_COEF => ROM20_DATA13_SIG,
    PE24_COEF => ROM20_DATA14_SIG,
    PE30_COEF => ROM20_DATA15_SIG,
    PE31_COEF => ROM20_DATA16_SIG,
    PE32_COEF => ROM20_DATA17_SIG,
    PE33_COEF => ROM20_DATA18_SIG,
    PE34_COEF => ROM20_DATA19_SIG,
    PE40_COEF => ROM20_DATA20_SIG,
    PE41_COEF => ROM20_DATA21_SIG,
    PE42_COEF => ROM20_DATA22_SIG,
    PE43_COEF => ROM20_DATA23_SIG,
    PE44_COEF => ROM20_DATA24_SIG,
    BIAS      => ROM20_DATA25_SIG,
    DOUT      => DOUT20_SIG
);

DSP_BLOCK21_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM21_DATA0_SIG,
    PE01_COEF => ROM21_DATA1_SIG,
    PE02_COEF => ROM21_DATA2_SIG,
    PE03_COEF => ROM21_DATA3_SIG,
    PE04_COEF => ROM21_DATA4_SIG,
    PE10_COEF => ROM21_DATA5_SIG,
    PE11_COEF => ROM21_DATA6_SIG,
    PE12_COEF => ROM21_DATA7_SIG,
    PE13_COEF => ROM21_DATA8_SIG,
    PE14_COEF => ROM21_DATA9_SIG,
    PE20_COEF => ROM21_DATA10_SIG,
    PE21_COEF => ROM21_DATA11_SIG,
    PE22_COEF => ROM21_DATA12_SIG,
    PE23_COEF => ROM21_DATA13_SIG,
    PE24_COEF => ROM21_DATA14_SIG,
    PE30_COEF => ROM21_DATA15_SIG,
    PE31_COEF => ROM21_DATA16_SIG,
    PE32_COEF => ROM21_DATA17_SIG,
    PE33_COEF => ROM21_DATA18_SIG,
    PE34_COEF => ROM21_DATA19_SIG,
    PE40_COEF => ROM21_DATA20_SIG,
    PE41_COEF => ROM21_DATA21_SIG,
    PE42_COEF => ROM21_DATA22_SIG,
    PE43_COEF => ROM21_DATA23_SIG,
    PE44_COEF => ROM21_DATA24_SIG,
    BIAS      => ROM21_DATA25_SIG,
    DOUT      => DOUT21_SIG
);

DSP_BLOCK22_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM22_DATA0_SIG,
    PE01_COEF => ROM22_DATA1_SIG,
    PE02_COEF => ROM22_DATA2_SIG,
    PE03_COEF => ROM22_DATA3_SIG,
    PE04_COEF => ROM22_DATA4_SIG,
    PE10_COEF => ROM22_DATA5_SIG,
    PE11_COEF => ROM22_DATA6_SIG,
    PE12_COEF => ROM22_DATA7_SIG,
    PE13_COEF => ROM22_DATA8_SIG,
    PE14_COEF => ROM22_DATA9_SIG,
    PE20_COEF => ROM22_DATA10_SIG,
    PE21_COEF => ROM22_DATA11_SIG,
    PE22_COEF => ROM22_DATA12_SIG,
    PE23_COEF => ROM22_DATA13_SIG,
    PE24_COEF => ROM22_DATA14_SIG,
    PE30_COEF => ROM22_DATA15_SIG,
    PE31_COEF => ROM22_DATA16_SIG,
    PE32_COEF => ROM22_DATA17_SIG,
    PE33_COEF => ROM22_DATA18_SIG,
    PE34_COEF => ROM22_DATA19_SIG,
    PE40_COEF => ROM22_DATA20_SIG,
    PE41_COEF => ROM22_DATA21_SIG,
    PE42_COEF => ROM22_DATA22_SIG,
    PE43_COEF => ROM22_DATA23_SIG,
    PE44_COEF => ROM22_DATA24_SIG,
    BIAS      => ROM22_DATA25_SIG,
    DOUT      => DOUT22_SIG
);

DSP_BLOCK23_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM23_DATA0_SIG,
    PE01_COEF => ROM23_DATA1_SIG,
    PE02_COEF => ROM23_DATA2_SIG,
    PE03_COEF => ROM23_DATA3_SIG,
    PE04_COEF => ROM23_DATA4_SIG,
    PE10_COEF => ROM23_DATA5_SIG,
    PE11_COEF => ROM23_DATA6_SIG,
    PE12_COEF => ROM23_DATA7_SIG,
    PE13_COEF => ROM23_DATA8_SIG,
    PE14_COEF => ROM23_DATA9_SIG,
    PE20_COEF => ROM23_DATA10_SIG,
    PE21_COEF => ROM23_DATA11_SIG,
    PE22_COEF => ROM23_DATA12_SIG,
    PE23_COEF => ROM23_DATA13_SIG,
    PE24_COEF => ROM23_DATA14_SIG,
    PE30_COEF => ROM23_DATA15_SIG,
    PE31_COEF => ROM23_DATA16_SIG,
    PE32_COEF => ROM23_DATA17_SIG,
    PE33_COEF => ROM23_DATA18_SIG,
    PE34_COEF => ROM23_DATA19_SIG,
    PE40_COEF => ROM23_DATA20_SIG,
    PE41_COEF => ROM23_DATA21_SIG,
    PE42_COEF => ROM23_DATA22_SIG,
    PE43_COEF => ROM23_DATA23_SIG,
    PE44_COEF => ROM23_DATA24_SIG,
    BIAS      => ROM23_DATA25_SIG,
    DOUT      => DOUT23_SIG
);

DSP_BLOCK24_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM24_DATA0_SIG,
    PE01_COEF => ROM24_DATA1_SIG,
    PE02_COEF => ROM24_DATA2_SIG,
    PE03_COEF => ROM24_DATA3_SIG,
    PE04_COEF => ROM24_DATA4_SIG,
    PE10_COEF => ROM24_DATA5_SIG,
    PE11_COEF => ROM24_DATA6_SIG,
    PE12_COEF => ROM24_DATA7_SIG,
    PE13_COEF => ROM24_DATA8_SIG,
    PE14_COEF => ROM24_DATA9_SIG,
    PE20_COEF => ROM24_DATA10_SIG,
    PE21_COEF => ROM24_DATA11_SIG,
    PE22_COEF => ROM24_DATA12_SIG,
    PE23_COEF => ROM24_DATA13_SIG,
    PE24_COEF => ROM24_DATA14_SIG,
    PE30_COEF => ROM24_DATA15_SIG,
    PE31_COEF => ROM24_DATA16_SIG,
    PE32_COEF => ROM24_DATA17_SIG,
    PE33_COEF => ROM24_DATA18_SIG,
    PE34_COEF => ROM24_DATA19_SIG,
    PE40_COEF => ROM24_DATA20_SIG,
    PE41_COEF => ROM24_DATA21_SIG,
    PE42_COEF => ROM24_DATA22_SIG,
    PE43_COEF => ROM24_DATA23_SIG,
    PE44_COEF => ROM24_DATA24_SIG,
    BIAS      => ROM24_DATA25_SIG,
    DOUT      => DOUT24_SIG
);

DSP_BLOCK25_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM25_DATA0_SIG,
    PE01_COEF => ROM25_DATA1_SIG,
    PE02_COEF => ROM25_DATA2_SIG,
    PE03_COEF => ROM25_DATA3_SIG,
    PE04_COEF => ROM25_DATA4_SIG,
    PE10_COEF => ROM25_DATA5_SIG,
    PE11_COEF => ROM25_DATA6_SIG,
    PE12_COEF => ROM25_DATA7_SIG,
    PE13_COEF => ROM25_DATA8_SIG,
    PE14_COEF => ROM25_DATA9_SIG,
    PE20_COEF => ROM25_DATA10_SIG,
    PE21_COEF => ROM25_DATA11_SIG,
    PE22_COEF => ROM25_DATA12_SIG,
    PE23_COEF => ROM25_DATA13_SIG,
    PE24_COEF => ROM25_DATA14_SIG,
    PE30_COEF => ROM25_DATA15_SIG,
    PE31_COEF => ROM25_DATA16_SIG,
    PE32_COEF => ROM25_DATA17_SIG,
    PE33_COEF => ROM25_DATA18_SIG,
    PE34_COEF => ROM25_DATA19_SIG,
    PE40_COEF => ROM25_DATA20_SIG,
    PE41_COEF => ROM25_DATA21_SIG,
    PE42_COEF => ROM25_DATA22_SIG,
    PE43_COEF => ROM25_DATA23_SIG,
    PE44_COEF => ROM25_DATA24_SIG,
    BIAS      => ROM25_DATA25_SIG,
    DOUT      => DOUT25_SIG
);

DSP_BLOCK26_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM26_DATA0_SIG,
    PE01_COEF => ROM26_DATA1_SIG,
    PE02_COEF => ROM26_DATA2_SIG,
    PE03_COEF => ROM26_DATA3_SIG,
    PE04_COEF => ROM26_DATA4_SIG,
    PE10_COEF => ROM26_DATA5_SIG,
    PE11_COEF => ROM26_DATA6_SIG,
    PE12_COEF => ROM26_DATA7_SIG,
    PE13_COEF => ROM26_DATA8_SIG,
    PE14_COEF => ROM26_DATA9_SIG,
    PE20_COEF => ROM26_DATA10_SIG,
    PE21_COEF => ROM26_DATA11_SIG,
    PE22_COEF => ROM26_DATA12_SIG,
    PE23_COEF => ROM26_DATA13_SIG,
    PE24_COEF => ROM26_DATA14_SIG,
    PE30_COEF => ROM26_DATA15_SIG,
    PE31_COEF => ROM26_DATA16_SIG,
    PE32_COEF => ROM26_DATA17_SIG,
    PE33_COEF => ROM26_DATA18_SIG,
    PE34_COEF => ROM26_DATA19_SIG,
    PE40_COEF => ROM26_DATA20_SIG,
    PE41_COEF => ROM26_DATA21_SIG,
    PE42_COEF => ROM26_DATA22_SIG,
    PE43_COEF => ROM26_DATA23_SIG,
    PE44_COEF => ROM26_DATA24_SIG,
    BIAS      => ROM26_DATA25_SIG,
    DOUT      => DOUT26_SIG
);

DSP_BLOCK27_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM27_DATA0_SIG,
    PE01_COEF => ROM27_DATA1_SIG,
    PE02_COEF => ROM27_DATA2_SIG,
    PE03_COEF => ROM27_DATA3_SIG,
    PE04_COEF => ROM27_DATA4_SIG,
    PE10_COEF => ROM27_DATA5_SIG,
    PE11_COEF => ROM27_DATA6_SIG,
    PE12_COEF => ROM27_DATA7_SIG,
    PE13_COEF => ROM27_DATA8_SIG,
    PE14_COEF => ROM27_DATA9_SIG,
    PE20_COEF => ROM27_DATA10_SIG,
    PE21_COEF => ROM27_DATA11_SIG,
    PE22_COEF => ROM27_DATA12_SIG,
    PE23_COEF => ROM27_DATA13_SIG,
    PE24_COEF => ROM27_DATA14_SIG,
    PE30_COEF => ROM27_DATA15_SIG,
    PE31_COEF => ROM27_DATA16_SIG,
    PE32_COEF => ROM27_DATA17_SIG,
    PE33_COEF => ROM27_DATA18_SIG,
    PE34_COEF => ROM27_DATA19_SIG,
    PE40_COEF => ROM27_DATA20_SIG,
    PE41_COEF => ROM27_DATA21_SIG,
    PE42_COEF => ROM27_DATA22_SIG,
    PE43_COEF => ROM27_DATA23_SIG,
    PE44_COEF => ROM27_DATA24_SIG,
    BIAS      => ROM27_DATA25_SIG,
    DOUT      => DOUT27_SIG
);

DSP_BLOCK28_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM28_DATA0_SIG,
    PE01_COEF => ROM28_DATA1_SIG,
    PE02_COEF => ROM28_DATA2_SIG,
    PE03_COEF => ROM28_DATA3_SIG,
    PE04_COEF => ROM28_DATA4_SIG,
    PE10_COEF => ROM28_DATA5_SIG,
    PE11_COEF => ROM28_DATA6_SIG,
    PE12_COEF => ROM28_DATA7_SIG,
    PE13_COEF => ROM28_DATA8_SIG,
    PE14_COEF => ROM28_DATA9_SIG,
    PE20_COEF => ROM28_DATA10_SIG,
    PE21_COEF => ROM28_DATA11_SIG,
    PE22_COEF => ROM28_DATA12_SIG,
    PE23_COEF => ROM28_DATA13_SIG,
    PE24_COEF => ROM28_DATA14_SIG,
    PE30_COEF => ROM28_DATA15_SIG,
    PE31_COEF => ROM28_DATA16_SIG,
    PE32_COEF => ROM28_DATA17_SIG,
    PE33_COEF => ROM28_DATA18_SIG,
    PE34_COEF => ROM28_DATA19_SIG,
    PE40_COEF => ROM28_DATA20_SIG,
    PE41_COEF => ROM28_DATA21_SIG,
    PE42_COEF => ROM28_DATA22_SIG,
    PE43_COEF => ROM28_DATA23_SIG,
    PE44_COEF => ROM28_DATA24_SIG,
    BIAS      => ROM28_DATA25_SIG,
    DOUT      => DOUT28_SIG
);

DSP_BLOCK29_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM29_DATA0_SIG,
    PE01_COEF => ROM29_DATA1_SIG,
    PE02_COEF => ROM29_DATA2_SIG,
    PE03_COEF => ROM29_DATA3_SIG,
    PE04_COEF => ROM29_DATA4_SIG,
    PE10_COEF => ROM29_DATA5_SIG,
    PE11_COEF => ROM29_DATA6_SIG,
    PE12_COEF => ROM29_DATA7_SIG,
    PE13_COEF => ROM29_DATA8_SIG,
    PE14_COEF => ROM29_DATA9_SIG,
    PE20_COEF => ROM29_DATA10_SIG,
    PE21_COEF => ROM29_DATA11_SIG,
    PE22_COEF => ROM29_DATA12_SIG,
    PE23_COEF => ROM29_DATA13_SIG,
    PE24_COEF => ROM29_DATA14_SIG,
    PE30_COEF => ROM29_DATA15_SIG,
    PE31_COEF => ROM29_DATA16_SIG,
    PE32_COEF => ROM29_DATA17_SIG,
    PE33_COEF => ROM29_DATA18_SIG,
    PE34_COEF => ROM29_DATA19_SIG,
    PE40_COEF => ROM29_DATA20_SIG,
    PE41_COEF => ROM29_DATA21_SIG,
    PE42_COEF => ROM29_DATA22_SIG,
    PE43_COEF => ROM29_DATA23_SIG,
    PE44_COEF => ROM29_DATA24_SIG,
    BIAS      => ROM29_DATA25_SIG,
    DOUT      => DOUT29_SIG
);

DSP_BLOCK30_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM30_DATA0_SIG,
    PE01_COEF => ROM30_DATA1_SIG,
    PE02_COEF => ROM30_DATA2_SIG,
    PE03_COEF => ROM30_DATA3_SIG,
    PE04_COEF => ROM30_DATA4_SIG,
    PE10_COEF => ROM30_DATA5_SIG,
    PE11_COEF => ROM30_DATA6_SIG,
    PE12_COEF => ROM30_DATA7_SIG,
    PE13_COEF => ROM30_DATA8_SIG,
    PE14_COEF => ROM30_DATA9_SIG,
    PE20_COEF => ROM30_DATA10_SIG,
    PE21_COEF => ROM30_DATA11_SIG,
    PE22_COEF => ROM30_DATA12_SIG,
    PE23_COEF => ROM30_DATA13_SIG,
    PE24_COEF => ROM30_DATA14_SIG,
    PE30_COEF => ROM30_DATA15_SIG,
    PE31_COEF => ROM30_DATA16_SIG,
    PE32_COEF => ROM30_DATA17_SIG,
    PE33_COEF => ROM30_DATA18_SIG,
    PE34_COEF => ROM30_DATA19_SIG,
    PE40_COEF => ROM30_DATA20_SIG,
    PE41_COEF => ROM30_DATA21_SIG,
    PE42_COEF => ROM30_DATA22_SIG,
    PE43_COEF => ROM30_DATA23_SIG,
    PE44_COEF => ROM30_DATA24_SIG,
    BIAS      => ROM30_DATA25_SIG,
    DOUT      => DOUT30_SIG
);

DSP_BLOCK31_INST: DSP_BLOCK
Generic map( PIXEL_SIZE => 16,
             POWER => 5)
Port map(
    CLK       => CLK,
    RESET     => RESET,
    DIN0      => DIN0_SIG,
    DIN1      => DIN1_SIG,
    DIN2      => DIN2_SIG,
    DIN3      => DIN3_SIG,
    DIN4      => DIN4_SIG,
    PE00_COEF => ROM31_DATA0_SIG,
    PE01_COEF => ROM31_DATA1_SIG,
    PE02_COEF => ROM31_DATA2_SIG,
    PE03_COEF => ROM31_DATA3_SIG,
    PE04_COEF => ROM31_DATA4_SIG,
    PE10_COEF => ROM31_DATA5_SIG,
    PE11_COEF => ROM31_DATA6_SIG,
    PE12_COEF => ROM31_DATA7_SIG,
    PE13_COEF => ROM31_DATA8_SIG,
    PE14_COEF => ROM31_DATA9_SIG,
    PE20_COEF => ROM31_DATA10_SIG,
    PE21_COEF => ROM31_DATA11_SIG,
    PE22_COEF => ROM31_DATA12_SIG,
    PE23_COEF => ROM31_DATA13_SIG,
    PE24_COEF => ROM31_DATA14_SIG,
    PE30_COEF => ROM31_DATA15_SIG,
    PE31_COEF => ROM31_DATA16_SIG,
    PE32_COEF => ROM31_DATA17_SIG,
    PE33_COEF => ROM31_DATA18_SIG,
    PE34_COEF => ROM31_DATA19_SIG,
    PE40_COEF => ROM31_DATA20_SIG,
    PE41_COEF => ROM31_DATA21_SIG,
    PE42_COEF => ROM31_DATA22_SIG,
    PE43_COEF => ROM31_DATA23_SIG,
    PE44_COEF => ROM31_DATA24_SIG,
    BIAS      => ROM31_DATA25_SIG,
    DOUT      => DOUT31_SIG
);

ROM0_INST: ROM0
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM0_DATA0_SIG,
    DATA1  => ROM0_DATA1_SIG,
    DATA2  => ROM0_DATA2_SIG,
    DATA3  => ROM0_DATA3_SIG,
    DATA4  => ROM0_DATA4_SIG,
    DATA5  => ROM0_DATA5_SIG,
    DATA6  => ROM0_DATA6_SIG,
    DATA7  => ROM0_DATA7_SIG,
    DATA8  => ROM0_DATA8_SIG,
    DATA9  => ROM0_DATA9_SIG,
    DATA10 => ROM0_DATA10_SIG,
    DATA11 => ROM0_DATA11_SIG,
    DATA12 => ROM0_DATA12_SIG,
    DATA13 => ROM0_DATA13_SIG,
    DATA14 => ROM0_DATA14_SIG,
    DATA15 => ROM0_DATA15_SIG,
    DATA16 => ROM0_DATA16_SIG,
    DATA17 => ROM0_DATA17_SIG,
    DATA18 => ROM0_DATA18_SIG,
    DATA19 => ROM0_DATA19_SIG,
    DATA20 => ROM0_DATA20_SIG,
    DATA21 => ROM0_DATA21_SIG,
    DATA22 => ROM0_DATA22_SIG,
    DATA23 => ROM0_DATA23_SIG,
    DATA24 => ROM0_DATA24_SIG,
    DATA25 => ROM0_DATA25_SIG
);

ROM1_INST: ROM1
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM1_DATA0_SIG,
    DATA1  => ROM1_DATA1_SIG,
    DATA2  => ROM1_DATA2_SIG,
    DATA3  => ROM1_DATA3_SIG,
    DATA4  => ROM1_DATA4_SIG,
    DATA5  => ROM1_DATA5_SIG,
    DATA6  => ROM1_DATA6_SIG,
    DATA7  => ROM1_DATA7_SIG,
    DATA8  => ROM1_DATA8_SIG,
    DATA9  => ROM1_DATA9_SIG,
    DATA10 => ROM1_DATA10_SIG,
    DATA11 => ROM1_DATA11_SIG,
    DATA12 => ROM1_DATA12_SIG,
    DATA13 => ROM1_DATA13_SIG,
    DATA14 => ROM1_DATA14_SIG,
    DATA15 => ROM1_DATA15_SIG,
    DATA16 => ROM1_DATA16_SIG,
    DATA17 => ROM1_DATA17_SIG,
    DATA18 => ROM1_DATA18_SIG,
    DATA19 => ROM1_DATA19_SIG,
    DATA20 => ROM1_DATA20_SIG,
    DATA21 => ROM1_DATA21_SIG,
    DATA22 => ROM1_DATA22_SIG,
    DATA23 => ROM1_DATA23_SIG,
    DATA24 => ROM1_DATA24_SIG,
    DATA25 => ROM1_DATA25_SIG
);

ROM2_INST: ROM2
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM2_DATA0_SIG,
    DATA1  => ROM2_DATA1_SIG,
    DATA2  => ROM2_DATA2_SIG,
    DATA3  => ROM2_DATA3_SIG,
    DATA4  => ROM2_DATA4_SIG,
    DATA5  => ROM2_DATA5_SIG,
    DATA6  => ROM2_DATA6_SIG,
    DATA7  => ROM2_DATA7_SIG,
    DATA8  => ROM2_DATA8_SIG,
    DATA9  => ROM2_DATA9_SIG,
    DATA10 => ROM2_DATA10_SIG,
    DATA11 => ROM2_DATA11_SIG,
    DATA12 => ROM2_DATA12_SIG,
    DATA13 => ROM2_DATA13_SIG,
    DATA14 => ROM2_DATA14_SIG,
    DATA15 => ROM2_DATA15_SIG,
    DATA16 => ROM2_DATA16_SIG,
    DATA17 => ROM2_DATA17_SIG,
    DATA18 => ROM2_DATA18_SIG,
    DATA19 => ROM2_DATA19_SIG,
    DATA20 => ROM2_DATA20_SIG,
    DATA21 => ROM2_DATA21_SIG,
    DATA22 => ROM2_DATA22_SIG,
    DATA23 => ROM2_DATA23_SIG,
    DATA24 => ROM2_DATA24_SIG,
    DATA25 => ROM2_DATA25_SIG
);

ROM3_INST: ROM3
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM3_DATA0_SIG,
    DATA1  => ROM3_DATA1_SIG,
    DATA2  => ROM3_DATA2_SIG,
    DATA3  => ROM3_DATA3_SIG,
    DATA4  => ROM3_DATA4_SIG,
    DATA5  => ROM3_DATA5_SIG,
    DATA6  => ROM3_DATA6_SIG,
    DATA7  => ROM3_DATA7_SIG,
    DATA8  => ROM3_DATA8_SIG,
    DATA9  => ROM3_DATA9_SIG,
    DATA10 => ROM3_DATA10_SIG,
    DATA11 => ROM3_DATA11_SIG,
    DATA12 => ROM3_DATA12_SIG,
    DATA13 => ROM3_DATA13_SIG,
    DATA14 => ROM3_DATA14_SIG,
    DATA15 => ROM3_DATA15_SIG,
    DATA16 => ROM3_DATA16_SIG,
    DATA17 => ROM3_DATA17_SIG,
    DATA18 => ROM3_DATA18_SIG,
    DATA19 => ROM3_DATA19_SIG,
    DATA20 => ROM3_DATA20_SIG,
    DATA21 => ROM3_DATA21_SIG,
    DATA22 => ROM3_DATA22_SIG,
    DATA23 => ROM3_DATA23_SIG,
    DATA24 => ROM3_DATA24_SIG,
    DATA25 => ROM3_DATA25_SIG
);

ROM4_INST: ROM4
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM4_DATA0_SIG,
    DATA1  => ROM4_DATA1_SIG,
    DATA2  => ROM4_DATA2_SIG,
    DATA3  => ROM4_DATA3_SIG,
    DATA4  => ROM4_DATA4_SIG,
    DATA5  => ROM4_DATA5_SIG,
    DATA6  => ROM4_DATA6_SIG,
    DATA7  => ROM4_DATA7_SIG,
    DATA8  => ROM4_DATA8_SIG,
    DATA9  => ROM4_DATA9_SIG,
    DATA10 => ROM4_DATA10_SIG,
    DATA11 => ROM4_DATA11_SIG,
    DATA12 => ROM4_DATA12_SIG,
    DATA13 => ROM4_DATA13_SIG,
    DATA14 => ROM4_DATA14_SIG,
    DATA15 => ROM4_DATA15_SIG,
    DATA16 => ROM4_DATA16_SIG,
    DATA17 => ROM4_DATA17_SIG,
    DATA18 => ROM4_DATA18_SIG,
    DATA19 => ROM4_DATA19_SIG,
    DATA20 => ROM4_DATA20_SIG,
    DATA21 => ROM4_DATA21_SIG,
    DATA22 => ROM4_DATA22_SIG,
    DATA23 => ROM4_DATA23_SIG,
    DATA24 => ROM4_DATA24_SIG,
    DATA25 => ROM4_DATA25_SIG
);

ROM5_INST: ROM5
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM5_DATA0_SIG,
    DATA1  => ROM5_DATA1_SIG,
    DATA2  => ROM5_DATA2_SIG,
    DATA3  => ROM5_DATA3_SIG,
    DATA4  => ROM5_DATA4_SIG,
    DATA5  => ROM5_DATA5_SIG,
    DATA6  => ROM5_DATA6_SIG,
    DATA7  => ROM5_DATA7_SIG,
    DATA8  => ROM5_DATA8_SIG,
    DATA9  => ROM5_DATA9_SIG,
    DATA10 => ROM5_DATA10_SIG,
    DATA11 => ROM5_DATA11_SIG,
    DATA12 => ROM5_DATA12_SIG,
    DATA13 => ROM5_DATA13_SIG,
    DATA14 => ROM5_DATA14_SIG,
    DATA15 => ROM5_DATA15_SIG,
    DATA16 => ROM5_DATA16_SIG,
    DATA17 => ROM5_DATA17_SIG,
    DATA18 => ROM5_DATA18_SIG,
    DATA19 => ROM5_DATA19_SIG,
    DATA20 => ROM5_DATA20_SIG,
    DATA21 => ROM5_DATA21_SIG,
    DATA22 => ROM5_DATA22_SIG,
    DATA23 => ROM5_DATA23_SIG,
    DATA24 => ROM5_DATA24_SIG,
    DATA25 => ROM5_DATA25_SIG
);

ROM6_INST: ROM6
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM6_DATA0_SIG,
    DATA1  => ROM6_DATA1_SIG,
    DATA2  => ROM6_DATA2_SIG,
    DATA3  => ROM6_DATA3_SIG,
    DATA4  => ROM6_DATA4_SIG,
    DATA5  => ROM6_DATA5_SIG,
    DATA6  => ROM6_DATA6_SIG,
    DATA7  => ROM6_DATA7_SIG,
    DATA8  => ROM6_DATA8_SIG,
    DATA9  => ROM6_DATA9_SIG,
    DATA10 => ROM6_DATA10_SIG,
    DATA11 => ROM6_DATA11_SIG,
    DATA12 => ROM6_DATA12_SIG,
    DATA13 => ROM6_DATA13_SIG,
    DATA14 => ROM6_DATA14_SIG,
    DATA15 => ROM6_DATA15_SIG,
    DATA16 => ROM6_DATA16_SIG,
    DATA17 => ROM6_DATA17_SIG,
    DATA18 => ROM6_DATA18_SIG,
    DATA19 => ROM6_DATA19_SIG,
    DATA20 => ROM6_DATA20_SIG,
    DATA21 => ROM6_DATA21_SIG,
    DATA22 => ROM6_DATA22_SIG,
    DATA23 => ROM6_DATA23_SIG,
    DATA24 => ROM6_DATA24_SIG,
    DATA25 => ROM6_DATA25_SIG
);

ROM7_INST: ROM7
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM7_DATA0_SIG,
    DATA1  => ROM7_DATA1_SIG,
    DATA2  => ROM7_DATA2_SIG,
    DATA3  => ROM7_DATA3_SIG,
    DATA4  => ROM7_DATA4_SIG,
    DATA5  => ROM7_DATA5_SIG,
    DATA6  => ROM7_DATA6_SIG,
    DATA7  => ROM7_DATA7_SIG,
    DATA8  => ROM7_DATA8_SIG,
    DATA9  => ROM7_DATA9_SIG,
    DATA10 => ROM7_DATA10_SIG,
    DATA11 => ROM7_DATA11_SIG,
    DATA12 => ROM7_DATA12_SIG,
    DATA13 => ROM7_DATA13_SIG,
    DATA14 => ROM7_DATA14_SIG,
    DATA15 => ROM7_DATA15_SIG,
    DATA16 => ROM7_DATA16_SIG,
    DATA17 => ROM7_DATA17_SIG,
    DATA18 => ROM7_DATA18_SIG,
    DATA19 => ROM7_DATA19_SIG,
    DATA20 => ROM7_DATA20_SIG,
    DATA21 => ROM7_DATA21_SIG,
    DATA22 => ROM7_DATA22_SIG,
    DATA23 => ROM7_DATA23_SIG,
    DATA24 => ROM7_DATA24_SIG,
    DATA25 => ROM7_DATA25_SIG
);

ROM8_INST: ROM8
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM8_DATA0_SIG,
    DATA1  => ROM8_DATA1_SIG,
    DATA2  => ROM8_DATA2_SIG,
    DATA3  => ROM8_DATA3_SIG,
    DATA4  => ROM8_DATA4_SIG,
    DATA5  => ROM8_DATA5_SIG,
    DATA6  => ROM8_DATA6_SIG,
    DATA7  => ROM8_DATA7_SIG,
    DATA8  => ROM8_DATA8_SIG,
    DATA9  => ROM8_DATA9_SIG,
    DATA10 => ROM8_DATA10_SIG,
    DATA11 => ROM8_DATA11_SIG,
    DATA12 => ROM8_DATA12_SIG,
    DATA13 => ROM8_DATA13_SIG,
    DATA14 => ROM8_DATA14_SIG,
    DATA15 => ROM8_DATA15_SIG,
    DATA16 => ROM8_DATA16_SIG,
    DATA17 => ROM8_DATA17_SIG,
    DATA18 => ROM8_DATA18_SIG,
    DATA19 => ROM8_DATA19_SIG,
    DATA20 => ROM8_DATA20_SIG,
    DATA21 => ROM8_DATA21_SIG,
    DATA22 => ROM8_DATA22_SIG,
    DATA23 => ROM8_DATA23_SIG,
    DATA24 => ROM8_DATA24_SIG,
    DATA25 => ROM8_DATA25_SIG
);

ROM9_INST: ROM9
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM9_DATA0_SIG,
    DATA1  => ROM9_DATA1_SIG,
    DATA2  => ROM9_DATA2_SIG,
    DATA3  => ROM9_DATA3_SIG,
    DATA4  => ROM9_DATA4_SIG,
    DATA5  => ROM9_DATA5_SIG,
    DATA6  => ROM9_DATA6_SIG,
    DATA7  => ROM9_DATA7_SIG,
    DATA8  => ROM9_DATA8_SIG,
    DATA9  => ROM9_DATA9_SIG,
    DATA10 => ROM9_DATA10_SIG,
    DATA11 => ROM9_DATA11_SIG,
    DATA12 => ROM9_DATA12_SIG,
    DATA13 => ROM9_DATA13_SIG,
    DATA14 => ROM9_DATA14_SIG,
    DATA15 => ROM9_DATA15_SIG,
    DATA16 => ROM9_DATA16_SIG,
    DATA17 => ROM9_DATA17_SIG,
    DATA18 => ROM9_DATA18_SIG,
    DATA19 => ROM9_DATA19_SIG,
    DATA20 => ROM9_DATA20_SIG,
    DATA21 => ROM9_DATA21_SIG,
    DATA22 => ROM9_DATA22_SIG,
    DATA23 => ROM9_DATA23_SIG,
    DATA24 => ROM9_DATA24_SIG,
    DATA25 => ROM9_DATA25_SIG
);

ROM10_INST: ROM10
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM10_DATA0_SIG,
    DATA1  => ROM10_DATA1_SIG,
    DATA2  => ROM10_DATA2_SIG,
    DATA3  => ROM10_DATA3_SIG,
    DATA4  => ROM10_DATA4_SIG,
    DATA5  => ROM10_DATA5_SIG,
    DATA6  => ROM10_DATA6_SIG,
    DATA7  => ROM10_DATA7_SIG,
    DATA8  => ROM10_DATA8_SIG,
    DATA9  => ROM10_DATA9_SIG,
    DATA10 => ROM10_DATA10_SIG,
    DATA11 => ROM10_DATA11_SIG,
    DATA12 => ROM10_DATA12_SIG,
    DATA13 => ROM10_DATA13_SIG,
    DATA14 => ROM10_DATA14_SIG,
    DATA15 => ROM10_DATA15_SIG,
    DATA16 => ROM10_DATA16_SIG,
    DATA17 => ROM10_DATA17_SIG,
    DATA18 => ROM10_DATA18_SIG,
    DATA19 => ROM10_DATA19_SIG,
    DATA20 => ROM10_DATA20_SIG,
    DATA21 => ROM10_DATA21_SIG,
    DATA22 => ROM10_DATA22_SIG,
    DATA23 => ROM10_DATA23_SIG,
    DATA24 => ROM10_DATA24_SIG,
    DATA25 => ROM10_DATA25_SIG
);

ROM11_INST: ROM11
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM11_DATA0_SIG,
    DATA1  => ROM11_DATA1_SIG,
    DATA2  => ROM11_DATA2_SIG,
    DATA3  => ROM11_DATA3_SIG,
    DATA4  => ROM11_DATA4_SIG,
    DATA5  => ROM11_DATA5_SIG,
    DATA6  => ROM11_DATA6_SIG,
    DATA7  => ROM11_DATA7_SIG,
    DATA8  => ROM11_DATA8_SIG,
    DATA9  => ROM11_DATA9_SIG,
    DATA10 => ROM11_DATA10_SIG,
    DATA11 => ROM11_DATA11_SIG,
    DATA12 => ROM11_DATA12_SIG,
    DATA13 => ROM11_DATA13_SIG,
    DATA14 => ROM11_DATA14_SIG,
    DATA15 => ROM11_DATA15_SIG,
    DATA16 => ROM11_DATA16_SIG,
    DATA17 => ROM11_DATA17_SIG,
    DATA18 => ROM11_DATA18_SIG,
    DATA19 => ROM11_DATA19_SIG,
    DATA20 => ROM11_DATA20_SIG,
    DATA21 => ROM11_DATA21_SIG,
    DATA22 => ROM11_DATA22_SIG,
    DATA23 => ROM11_DATA23_SIG,
    DATA24 => ROM11_DATA24_SIG,
    DATA25 => ROM11_DATA25_SIG
);

ROM12_INST: ROM12
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM12_DATA0_SIG,
    DATA1  => ROM12_DATA1_SIG,
    DATA2  => ROM12_DATA2_SIG,
    DATA3  => ROM12_DATA3_SIG,
    DATA4  => ROM12_DATA4_SIG,
    DATA5  => ROM12_DATA5_SIG,
    DATA6  => ROM12_DATA6_SIG,
    DATA7  => ROM12_DATA7_SIG,
    DATA8  => ROM12_DATA8_SIG,
    DATA9  => ROM12_DATA9_SIG,
    DATA10 => ROM12_DATA10_SIG,
    DATA11 => ROM12_DATA11_SIG,
    DATA12 => ROM12_DATA12_SIG,
    DATA13 => ROM12_DATA13_SIG,
    DATA14 => ROM12_DATA14_SIG,
    DATA15 => ROM12_DATA15_SIG,
    DATA16 => ROM12_DATA16_SIG,
    DATA17 => ROM12_DATA17_SIG,
    DATA18 => ROM12_DATA18_SIG,
    DATA19 => ROM12_DATA19_SIG,
    DATA20 => ROM12_DATA20_SIG,
    DATA21 => ROM12_DATA21_SIG,
    DATA22 => ROM12_DATA22_SIG,
    DATA23 => ROM12_DATA23_SIG,
    DATA24 => ROM12_DATA24_SIG,
    DATA25 => ROM12_DATA25_SIG
);

ROM13_INST: ROM13
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM13_DATA0_SIG,
    DATA1  => ROM13_DATA1_SIG,
    DATA2  => ROM13_DATA2_SIG,
    DATA3  => ROM13_DATA3_SIG,
    DATA4  => ROM13_DATA4_SIG,
    DATA5  => ROM13_DATA5_SIG,
    DATA6  => ROM13_DATA6_SIG,
    DATA7  => ROM13_DATA7_SIG,
    DATA8  => ROM13_DATA8_SIG,
    DATA9  => ROM13_DATA9_SIG,
    DATA10 => ROM13_DATA10_SIG,
    DATA11 => ROM13_DATA11_SIG,
    DATA12 => ROM13_DATA12_SIG,
    DATA13 => ROM13_DATA13_SIG,
    DATA14 => ROM13_DATA14_SIG,
    DATA15 => ROM13_DATA15_SIG,
    DATA16 => ROM13_DATA16_SIG,
    DATA17 => ROM13_DATA17_SIG,
    DATA18 => ROM13_DATA18_SIG,
    DATA19 => ROM13_DATA19_SIG,
    DATA20 => ROM13_DATA20_SIG,
    DATA21 => ROM13_DATA21_SIG,
    DATA22 => ROM13_DATA22_SIG,
    DATA23 => ROM13_DATA23_SIG,
    DATA24 => ROM13_DATA24_SIG,
    DATA25 => ROM13_DATA25_SIG
);

ROM14_INST: ROM14
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM14_DATA0_SIG,
    DATA1  => ROM14_DATA1_SIG,
    DATA2  => ROM14_DATA2_SIG,
    DATA3  => ROM14_DATA3_SIG,
    DATA4  => ROM14_DATA4_SIG,
    DATA5  => ROM14_DATA5_SIG,
    DATA6  => ROM14_DATA6_SIG,
    DATA7  => ROM14_DATA7_SIG,
    DATA8  => ROM14_DATA8_SIG,
    DATA9  => ROM14_DATA9_SIG,
    DATA10 => ROM14_DATA10_SIG,
    DATA11 => ROM14_DATA11_SIG,
    DATA12 => ROM14_DATA12_SIG,
    DATA13 => ROM14_DATA13_SIG,
    DATA14 => ROM14_DATA14_SIG,
    DATA15 => ROM14_DATA15_SIG,
    DATA16 => ROM14_DATA16_SIG,
    DATA17 => ROM14_DATA17_SIG,
    DATA18 => ROM14_DATA18_SIG,
    DATA19 => ROM14_DATA19_SIG,
    DATA20 => ROM14_DATA20_SIG,
    DATA21 => ROM14_DATA21_SIG,
    DATA22 => ROM14_DATA22_SIG,
    DATA23 => ROM14_DATA23_SIG,
    DATA24 => ROM14_DATA24_SIG,
    DATA25 => ROM14_DATA25_SIG
);

ROM15_INST: ROM15
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM15_DATA0_SIG,
    DATA1  => ROM15_DATA1_SIG,
    DATA2  => ROM15_DATA2_SIG,
    DATA3  => ROM15_DATA3_SIG,
    DATA4  => ROM15_DATA4_SIG,
    DATA5  => ROM15_DATA5_SIG,
    DATA6  => ROM15_DATA6_SIG,
    DATA7  => ROM15_DATA7_SIG,
    DATA8  => ROM15_DATA8_SIG,
    DATA9  => ROM15_DATA9_SIG,
    DATA10 => ROM15_DATA10_SIG,
    DATA11 => ROM15_DATA11_SIG,
    DATA12 => ROM15_DATA12_SIG,
    DATA13 => ROM15_DATA13_SIG,
    DATA14 => ROM15_DATA14_SIG,
    DATA15 => ROM15_DATA15_SIG,
    DATA16 => ROM15_DATA16_SIG,
    DATA17 => ROM15_DATA17_SIG,
    DATA18 => ROM15_DATA18_SIG,
    DATA19 => ROM15_DATA19_SIG,
    DATA20 => ROM15_DATA20_SIG,
    DATA21 => ROM15_DATA21_SIG,
    DATA22 => ROM15_DATA22_SIG,
    DATA23 => ROM15_DATA23_SIG,
    DATA24 => ROM15_DATA24_SIG,
    DATA25 => ROM15_DATA25_SIG
);

ROM16_INST: ROM16
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM16_DATA0_SIG,
    DATA1  => ROM16_DATA1_SIG,
    DATA2  => ROM16_DATA2_SIG,
    DATA3  => ROM16_DATA3_SIG,
    DATA4  => ROM16_DATA4_SIG,
    DATA5  => ROM16_DATA5_SIG,
    DATA6  => ROM16_DATA6_SIG,
    DATA7  => ROM16_DATA7_SIG,
    DATA8  => ROM16_DATA8_SIG,
    DATA9  => ROM16_DATA9_SIG,
    DATA10 => ROM16_DATA10_SIG,
    DATA11 => ROM16_DATA11_SIG,
    DATA12 => ROM16_DATA12_SIG,
    DATA13 => ROM16_DATA13_SIG,
    DATA14 => ROM16_DATA14_SIG,
    DATA15 => ROM16_DATA15_SIG,
    DATA16 => ROM16_DATA16_SIG,
    DATA17 => ROM16_DATA17_SIG,
    DATA18 => ROM16_DATA18_SIG,
    DATA19 => ROM16_DATA19_SIG,
    DATA20 => ROM16_DATA20_SIG,
    DATA21 => ROM16_DATA21_SIG,
    DATA22 => ROM16_DATA22_SIG,
    DATA23 => ROM16_DATA23_SIG,
    DATA24 => ROM16_DATA24_SIG,
    DATA25 => ROM16_DATA25_SIG
);

ROM17_INST: ROM17
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM17_DATA0_SIG,
    DATA1  => ROM17_DATA1_SIG,
    DATA2  => ROM17_DATA2_SIG,
    DATA3  => ROM17_DATA3_SIG,
    DATA4  => ROM17_DATA4_SIG,
    DATA5  => ROM17_DATA5_SIG,
    DATA6  => ROM17_DATA6_SIG,
    DATA7  => ROM17_DATA7_SIG,
    DATA8  => ROM17_DATA8_SIG,
    DATA9  => ROM17_DATA9_SIG,
    DATA10 => ROM17_DATA10_SIG,
    DATA11 => ROM17_DATA11_SIG,
    DATA12 => ROM17_DATA12_SIG,
    DATA13 => ROM17_DATA13_SIG,
    DATA14 => ROM17_DATA14_SIG,
    DATA15 => ROM17_DATA15_SIG,
    DATA16 => ROM17_DATA16_SIG,
    DATA17 => ROM17_DATA17_SIG,
    DATA18 => ROM17_DATA18_SIG,
    DATA19 => ROM17_DATA19_SIG,
    DATA20 => ROM17_DATA20_SIG,
    DATA21 => ROM17_DATA21_SIG,
    DATA22 => ROM17_DATA22_SIG,
    DATA23 => ROM17_DATA23_SIG,
    DATA24 => ROM17_DATA24_SIG,
    DATA25 => ROM17_DATA25_SIG
);

ROM18_INST: ROM18
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM18_DATA0_SIG,
    DATA1  => ROM18_DATA1_SIG,
    DATA2  => ROM18_DATA2_SIG,
    DATA3  => ROM18_DATA3_SIG,
    DATA4  => ROM18_DATA4_SIG,
    DATA5  => ROM18_DATA5_SIG,
    DATA6  => ROM18_DATA6_SIG,
    DATA7  => ROM18_DATA7_SIG,
    DATA8  => ROM18_DATA8_SIG,
    DATA9  => ROM18_DATA9_SIG,
    DATA10 => ROM18_DATA10_SIG,
    DATA11 => ROM18_DATA11_SIG,
    DATA12 => ROM18_DATA12_SIG,
    DATA13 => ROM18_DATA13_SIG,
    DATA14 => ROM18_DATA14_SIG,
    DATA15 => ROM18_DATA15_SIG,
    DATA16 => ROM18_DATA16_SIG,
    DATA17 => ROM18_DATA17_SIG,
    DATA18 => ROM18_DATA18_SIG,
    DATA19 => ROM18_DATA19_SIG,
    DATA20 => ROM18_DATA20_SIG,
    DATA21 => ROM18_DATA21_SIG,
    DATA22 => ROM18_DATA22_SIG,
    DATA23 => ROM18_DATA23_SIG,
    DATA24 => ROM18_DATA24_SIG,
    DATA25 => ROM18_DATA25_SIG
);

ROM19_INST: ROM19
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM19_DATA0_SIG,
    DATA1  => ROM19_DATA1_SIG,
    DATA2  => ROM19_DATA2_SIG,
    DATA3  => ROM19_DATA3_SIG,
    DATA4  => ROM19_DATA4_SIG,
    DATA5  => ROM19_DATA5_SIG,
    DATA6  => ROM19_DATA6_SIG,
    DATA7  => ROM19_DATA7_SIG,
    DATA8  => ROM19_DATA8_SIG,
    DATA9  => ROM19_DATA9_SIG,
    DATA10 => ROM19_DATA10_SIG,
    DATA11 => ROM19_DATA11_SIG,
    DATA12 => ROM19_DATA12_SIG,
    DATA13 => ROM19_DATA13_SIG,
    DATA14 => ROM19_DATA14_SIG,
    DATA15 => ROM19_DATA15_SIG,
    DATA16 => ROM19_DATA16_SIG,
    DATA17 => ROM19_DATA17_SIG,
    DATA18 => ROM19_DATA18_SIG,
    DATA19 => ROM19_DATA19_SIG,
    DATA20 => ROM19_DATA20_SIG,
    DATA21 => ROM19_DATA21_SIG,
    DATA22 => ROM19_DATA22_SIG,
    DATA23 => ROM19_DATA23_SIG,
    DATA24 => ROM19_DATA24_SIG,
    DATA25 => ROM19_DATA25_SIG
);

ROM20_INST: ROM20
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM20_DATA0_SIG,
    DATA1  => ROM20_DATA1_SIG,
    DATA2  => ROM20_DATA2_SIG,
    DATA3  => ROM20_DATA3_SIG,
    DATA4  => ROM20_DATA4_SIG,
    DATA5  => ROM20_DATA5_SIG,
    DATA6  => ROM20_DATA6_SIG,
    DATA7  => ROM20_DATA7_SIG,
    DATA8  => ROM20_DATA8_SIG,
    DATA9  => ROM20_DATA9_SIG,
    DATA10 => ROM20_DATA10_SIG,
    DATA11 => ROM20_DATA11_SIG,
    DATA12 => ROM20_DATA12_SIG,
    DATA13 => ROM20_DATA13_SIG,
    DATA14 => ROM20_DATA14_SIG,
    DATA15 => ROM20_DATA15_SIG,
    DATA16 => ROM20_DATA16_SIG,
    DATA17 => ROM20_DATA17_SIG,
    DATA18 => ROM20_DATA18_SIG,
    DATA19 => ROM20_DATA19_SIG,
    DATA20 => ROM20_DATA20_SIG,
    DATA21 => ROM20_DATA21_SIG,
    DATA22 => ROM20_DATA22_SIG,
    DATA23 => ROM20_DATA23_SIG,
    DATA24 => ROM20_DATA24_SIG,
    DATA25 => ROM20_DATA25_SIG
);

ROM21_INST: ROM21
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM21_DATA0_SIG,
    DATA1  => ROM21_DATA1_SIG,
    DATA2  => ROM21_DATA2_SIG,
    DATA3  => ROM21_DATA3_SIG,
    DATA4  => ROM21_DATA4_SIG,
    DATA5  => ROM21_DATA5_SIG,
    DATA6  => ROM21_DATA6_SIG,
    DATA7  => ROM21_DATA7_SIG,
    DATA8  => ROM21_DATA8_SIG,
    DATA9  => ROM21_DATA9_SIG,
    DATA10 => ROM21_DATA10_SIG,
    DATA11 => ROM21_DATA11_SIG,
    DATA12 => ROM21_DATA12_SIG,
    DATA13 => ROM21_DATA13_SIG,
    DATA14 => ROM21_DATA14_SIG,
    DATA15 => ROM21_DATA15_SIG,
    DATA16 => ROM21_DATA16_SIG,
    DATA17 => ROM21_DATA17_SIG,
    DATA18 => ROM21_DATA18_SIG,
    DATA19 => ROM21_DATA19_SIG,
    DATA20 => ROM21_DATA20_SIG,
    DATA21 => ROM21_DATA21_SIG,
    DATA22 => ROM21_DATA22_SIG,
    DATA23 => ROM21_DATA23_SIG,
    DATA24 => ROM21_DATA24_SIG,
    DATA25 => ROM21_DATA25_SIG
);

ROM22_INST: ROM22
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM22_DATA0_SIG,
    DATA1  => ROM22_DATA1_SIG,
    DATA2  => ROM22_DATA2_SIG,
    DATA3  => ROM22_DATA3_SIG,
    DATA4  => ROM22_DATA4_SIG,
    DATA5  => ROM22_DATA5_SIG,
    DATA6  => ROM22_DATA6_SIG,
    DATA7  => ROM22_DATA7_SIG,
    DATA8  => ROM22_DATA8_SIG,
    DATA9  => ROM22_DATA9_SIG,
    DATA10 => ROM22_DATA10_SIG,
    DATA11 => ROM22_DATA11_SIG,
    DATA12 => ROM22_DATA12_SIG,
    DATA13 => ROM22_DATA13_SIG,
    DATA14 => ROM22_DATA14_SIG,
    DATA15 => ROM22_DATA15_SIG,
    DATA16 => ROM22_DATA16_SIG,
    DATA17 => ROM22_DATA17_SIG,
    DATA18 => ROM22_DATA18_SIG,
    DATA19 => ROM22_DATA19_SIG,
    DATA20 => ROM22_DATA20_SIG,
    DATA21 => ROM22_DATA21_SIG,
    DATA22 => ROM22_DATA22_SIG,
    DATA23 => ROM22_DATA23_SIG,
    DATA24 => ROM22_DATA24_SIG,
    DATA25 => ROM22_DATA25_SIG
);

ROM23_INST: ROM23
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM23_DATA0_SIG,
    DATA1  => ROM23_DATA1_SIG,
    DATA2  => ROM23_DATA2_SIG,
    DATA3  => ROM23_DATA3_SIG,
    DATA4  => ROM23_DATA4_SIG,
    DATA5  => ROM23_DATA5_SIG,
    DATA6  => ROM23_DATA6_SIG,
    DATA7  => ROM23_DATA7_SIG,
    DATA8  => ROM23_DATA8_SIG,
    DATA9  => ROM23_DATA9_SIG,
    DATA10 => ROM23_DATA10_SIG,
    DATA11 => ROM23_DATA11_SIG,
    DATA12 => ROM23_DATA12_SIG,
    DATA13 => ROM23_DATA13_SIG,
    DATA14 => ROM23_DATA14_SIG,
    DATA15 => ROM23_DATA15_SIG,
    DATA16 => ROM23_DATA16_SIG,
    DATA17 => ROM23_DATA17_SIG,
    DATA18 => ROM23_DATA18_SIG,
    DATA19 => ROM23_DATA19_SIG,
    DATA20 => ROM23_DATA20_SIG,
    DATA21 => ROM23_DATA21_SIG,
    DATA22 => ROM23_DATA22_SIG,
    DATA23 => ROM23_DATA23_SIG,
    DATA24 => ROM23_DATA24_SIG,
    DATA25 => ROM23_DATA25_SIG
);

ROM24_INST: ROM24
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM24_DATA0_SIG,
    DATA1  => ROM24_DATA1_SIG,
    DATA2  => ROM24_DATA2_SIG,
    DATA3  => ROM24_DATA3_SIG,
    DATA4  => ROM24_DATA4_SIG,
    DATA5  => ROM24_DATA5_SIG,
    DATA6  => ROM24_DATA6_SIG,
    DATA7  => ROM24_DATA7_SIG,
    DATA8  => ROM24_DATA8_SIG,
    DATA9  => ROM24_DATA9_SIG,
    DATA10 => ROM24_DATA10_SIG,
    DATA11 => ROM24_DATA11_SIG,
    DATA12 => ROM24_DATA12_SIG,
    DATA13 => ROM24_DATA13_SIG,
    DATA14 => ROM24_DATA14_SIG,
    DATA15 => ROM24_DATA15_SIG,
    DATA16 => ROM24_DATA16_SIG,
    DATA17 => ROM24_DATA17_SIG,
    DATA18 => ROM24_DATA18_SIG,
    DATA19 => ROM24_DATA19_SIG,
    DATA20 => ROM24_DATA20_SIG,
    DATA21 => ROM24_DATA21_SIG,
    DATA22 => ROM24_DATA22_SIG,
    DATA23 => ROM24_DATA23_SIG,
    DATA24 => ROM24_DATA24_SIG,
    DATA25 => ROM24_DATA25_SIG
);

ROM25_INST: ROM25
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM25_DATA0_SIG,
    DATA1  => ROM25_DATA1_SIG,
    DATA2  => ROM25_DATA2_SIG,
    DATA3  => ROM25_DATA3_SIG,
    DATA4  => ROM25_DATA4_SIG,
    DATA5  => ROM25_DATA5_SIG,
    DATA6  => ROM25_DATA6_SIG,
    DATA7  => ROM25_DATA7_SIG,
    DATA8  => ROM25_DATA8_SIG,
    DATA9  => ROM25_DATA9_SIG,
    DATA10 => ROM25_DATA10_SIG,
    DATA11 => ROM25_DATA11_SIG,
    DATA12 => ROM25_DATA12_SIG,
    DATA13 => ROM25_DATA13_SIG,
    DATA14 => ROM25_DATA14_SIG,
    DATA15 => ROM25_DATA15_SIG,
    DATA16 => ROM25_DATA16_SIG,
    DATA17 => ROM25_DATA17_SIG,
    DATA18 => ROM25_DATA18_SIG,
    DATA19 => ROM25_DATA19_SIG,
    DATA20 => ROM25_DATA20_SIG,
    DATA21 => ROM25_DATA21_SIG,
    DATA22 => ROM25_DATA22_SIG,
    DATA23 => ROM25_DATA23_SIG,
    DATA24 => ROM25_DATA24_SIG,
    DATA25 => ROM25_DATA25_SIG
);

ROM26_INST: ROM26
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM26_DATA0_SIG,
    DATA1  => ROM26_DATA1_SIG,
    DATA2  => ROM26_DATA2_SIG,
    DATA3  => ROM26_DATA3_SIG,
    DATA4  => ROM26_DATA4_SIG,
    DATA5  => ROM26_DATA5_SIG,
    DATA6  => ROM26_DATA6_SIG,
    DATA7  => ROM26_DATA7_SIG,
    DATA8  => ROM26_DATA8_SIG,
    DATA9  => ROM26_DATA9_SIG,
    DATA10 => ROM26_DATA10_SIG,
    DATA11 => ROM26_DATA11_SIG,
    DATA12 => ROM26_DATA12_SIG,
    DATA13 => ROM26_DATA13_SIG,
    DATA14 => ROM26_DATA14_SIG,
    DATA15 => ROM26_DATA15_SIG,
    DATA16 => ROM26_DATA16_SIG,
    DATA17 => ROM26_DATA17_SIG,
    DATA18 => ROM26_DATA18_SIG,
    DATA19 => ROM26_DATA19_SIG,
    DATA20 => ROM26_DATA20_SIG,
    DATA21 => ROM26_DATA21_SIG,
    DATA22 => ROM26_DATA22_SIG,
    DATA23 => ROM26_DATA23_SIG,
    DATA24 => ROM26_DATA24_SIG,
    DATA25 => ROM26_DATA25_SIG
);

ROM27_INST: ROM27
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM27_DATA0_SIG,
    DATA1  => ROM27_DATA1_SIG,
    DATA2  => ROM27_DATA2_SIG,
    DATA3  => ROM27_DATA3_SIG,
    DATA4  => ROM27_DATA4_SIG,
    DATA5  => ROM27_DATA5_SIG,
    DATA6  => ROM27_DATA6_SIG,
    DATA7  => ROM27_DATA7_SIG,
    DATA8  => ROM27_DATA8_SIG,
    DATA9  => ROM27_DATA9_SIG,
    DATA10 => ROM27_DATA10_SIG,
    DATA11 => ROM27_DATA11_SIG,
    DATA12 => ROM27_DATA12_SIG,
    DATA13 => ROM27_DATA13_SIG,
    DATA14 => ROM27_DATA14_SIG,
    DATA15 => ROM27_DATA15_SIG,
    DATA16 => ROM27_DATA16_SIG,
    DATA17 => ROM27_DATA17_SIG,
    DATA18 => ROM27_DATA18_SIG,
    DATA19 => ROM27_DATA19_SIG,
    DATA20 => ROM27_DATA20_SIG,
    DATA21 => ROM27_DATA21_SIG,
    DATA22 => ROM27_DATA22_SIG,
    DATA23 => ROM27_DATA23_SIG,
    DATA24 => ROM27_DATA24_SIG,
    DATA25 => ROM27_DATA25_SIG
);

ROM28_INST: ROM28
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM28_DATA0_SIG,
    DATA1  => ROM28_DATA1_SIG,
    DATA2  => ROM28_DATA2_SIG,
    DATA3  => ROM28_DATA3_SIG,
    DATA4  => ROM28_DATA4_SIG,
    DATA5  => ROM28_DATA5_SIG,
    DATA6  => ROM28_DATA6_SIG,
    DATA7  => ROM28_DATA7_SIG,
    DATA8  => ROM28_DATA8_SIG,
    DATA9  => ROM28_DATA9_SIG,
    DATA10 => ROM28_DATA10_SIG,
    DATA11 => ROM28_DATA11_SIG,
    DATA12 => ROM28_DATA12_SIG,
    DATA13 => ROM28_DATA13_SIG,
    DATA14 => ROM28_DATA14_SIG,
    DATA15 => ROM28_DATA15_SIG,
    DATA16 => ROM28_DATA16_SIG,
    DATA17 => ROM28_DATA17_SIG,
    DATA18 => ROM28_DATA18_SIG,
    DATA19 => ROM28_DATA19_SIG,
    DATA20 => ROM28_DATA20_SIG,
    DATA21 => ROM28_DATA21_SIG,
    DATA22 => ROM28_DATA22_SIG,
    DATA23 => ROM28_DATA23_SIG,
    DATA24 => ROM28_DATA24_SIG,
    DATA25 => ROM28_DATA25_SIG
);

ROM29_INST: ROM29
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM29_DATA0_SIG,
    DATA1  => ROM29_DATA1_SIG,
    DATA2  => ROM29_DATA2_SIG,
    DATA3  => ROM29_DATA3_SIG,
    DATA4  => ROM29_DATA4_SIG,
    DATA5  => ROM29_DATA5_SIG,
    DATA6  => ROM29_DATA6_SIG,
    DATA7  => ROM29_DATA7_SIG,
    DATA8  => ROM29_DATA8_SIG,
    DATA9  => ROM29_DATA9_SIG,
    DATA10 => ROM29_DATA10_SIG,
    DATA11 => ROM29_DATA11_SIG,
    DATA12 => ROM29_DATA12_SIG,
    DATA13 => ROM29_DATA13_SIG,
    DATA14 => ROM29_DATA14_SIG,
    DATA15 => ROM29_DATA15_SIG,
    DATA16 => ROM29_DATA16_SIG,
    DATA17 => ROM29_DATA17_SIG,
    DATA18 => ROM29_DATA18_SIG,
    DATA19 => ROM29_DATA19_SIG,
    DATA20 => ROM29_DATA20_SIG,
    DATA21 => ROM29_DATA21_SIG,
    DATA22 => ROM29_DATA22_SIG,
    DATA23 => ROM29_DATA23_SIG,
    DATA24 => ROM29_DATA24_SIG,
    DATA25 => ROM29_DATA25_SIG
);

ROM30_INST: ROM30
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM30_DATA0_SIG,
    DATA1  => ROM30_DATA1_SIG,
    DATA2  => ROM30_DATA2_SIG,
    DATA3  => ROM30_DATA3_SIG,
    DATA4  => ROM30_DATA4_SIG,
    DATA5  => ROM30_DATA5_SIG,
    DATA6  => ROM30_DATA6_SIG,
    DATA7  => ROM30_DATA7_SIG,
    DATA8  => ROM30_DATA8_SIG,
    DATA9  => ROM30_DATA9_SIG,
    DATA10 => ROM30_DATA10_SIG,
    DATA11 => ROM30_DATA11_SIG,
    DATA12 => ROM30_DATA12_SIG,
    DATA13 => ROM30_DATA13_SIG,
    DATA14 => ROM30_DATA14_SIG,
    DATA15 => ROM30_DATA15_SIG,
    DATA16 => ROM30_DATA16_SIG,
    DATA17 => ROM30_DATA17_SIG,
    DATA18 => ROM30_DATA18_SIG,
    DATA19 => ROM30_DATA19_SIG,
    DATA20 => ROM30_DATA20_SIG,
    DATA21 => ROM30_DATA21_SIG,
    DATA22 => ROM30_DATA22_SIG,
    DATA23 => ROM30_DATA23_SIG,
    DATA24 => ROM30_DATA24_SIG,
    DATA25 => ROM30_DATA25_SIG
);

ROM31_INST: ROM31
Generic map( WIDTH => 16,
          POWER => 5) 
Port map( 
    ADDR0  => ADDR0_SIG,
    ADDR1  => ADDR1_SIG,
    ADDR2  => ADDR2_SIG,
    ADDR3  => ADDR3_SIG,
    ADDR4  => ADDR4_SIG,
    ADDR5  => ADDR5_SIG,
    ADDR6  => ADDR6_SIG,
    ADDR7  => ADDR7_SIG,
    ADDR8  => ADDR8_SIG,
    ADDR9  => ADDR9_SIG,
    ADDR10 => ADDR10_SIG,
    ADDR11 => ADDR11_SIG,
    ADDR12 => ADDR12_SIG,
    ADDR13 => ADDR13_SIG,
    ADDR14 => ADDR14_SIG,
    ADDR15 => ADDR15_SIG,
    ADDR16 => ADDR16_SIG,
    ADDR17 => ADDR17_SIG,
    ADDR18 => ADDR18_SIG,
    ADDR19 => ADDR19_SIG,
    ADDR20 => ADDR20_SIG,
    ADDR21 => ADDR21_SIG,
    ADDR22 => ADDR22_SIG,
    ADDR23 => ADDR23_SIG,
    ADDR24 => ADDR24_SIG,
    ADDR25 => ADDR25_SIG,
    DATA0  => ROM31_DATA0_SIG,
    DATA1  => ROM31_DATA1_SIG,
    DATA2  => ROM31_DATA2_SIG,
    DATA3  => ROM31_DATA3_SIG,
    DATA4  => ROM31_DATA4_SIG,
    DATA5  => ROM31_DATA5_SIG,
    DATA6  => ROM31_DATA6_SIG,
    DATA7  => ROM31_DATA7_SIG,
    DATA8  => ROM31_DATA8_SIG,
    DATA9  => ROM31_DATA9_SIG,
    DATA10 => ROM31_DATA10_SIG,
    DATA11 => ROM31_DATA11_SIG,
    DATA12 => ROM31_DATA12_SIG,
    DATA13 => ROM31_DATA13_SIG,
    DATA14 => ROM31_DATA14_SIG,
    DATA15 => ROM31_DATA15_SIG,
    DATA16 => ROM31_DATA16_SIG,
    DATA17 => ROM31_DATA17_SIG,
    DATA18 => ROM31_DATA18_SIG,
    DATA19 => ROM31_DATA19_SIG,
    DATA20 => ROM31_DATA20_SIG,
    DATA21 => ROM31_DATA21_SIG,
    DATA22 => ROM31_DATA22_SIG,
    DATA23 => ROM31_DATA23_SIG,
    DATA24 => ROM31_DATA24_SIG,
    DATA25 => ROM31_DATA25_SIG
);

DOUT0 <= DOUT0_SIG;
DOUT1 <= DOUT1_SIG;
DOUT2 <= DOUT2_SIG;
DOUT3 <= DOUT3_SIG;
DOUT4 <= DOUT4_SIG;
DOUT5 <= DOUT5_SIG;
DOUT6 <= DOUT6_SIG;
DOUT7 <= DOUT7_SIG;
DOUT8 <= DOUT8_SIG;
DOUT9 <= DOUT9_SIG;
DOUT10 <= DOUT10_SIG;
DOUT11 <= DOUT11_SIG;
DOUT12 <= DOUT12_SIG;
DOUT13 <= DOUT13_SIG;
DOUT14 <= DOUT14_SIG;
DOUT15 <= DOUT15_SIG;
DOUT16 <= DOUT16_SIG;
DOUT17 <= DOUT17_SIG;
DOUT18 <= DOUT18_SIG;
DOUT19 <= DOUT19_SIG;
DOUT20 <= DOUT20_SIG;
DOUT21 <= DOUT21_SIG;
DOUT22 <= DOUT22_SIG;
DOUT23 <= DOUT23_SIG;
DOUT24 <= DOUT24_SIG;
DOUT25 <= DOUT25_SIG;
DOUT26 <= DOUT26_SIG;
DOUT27 <= DOUT27_SIG;
DOUT28 <= DOUT28_SIG;
DOUT29 <= DOUT29_SIG;
DOUT30 <= DOUT30_SIG;
DOUT31 <= DOUT31_SIG;

end Structural;
